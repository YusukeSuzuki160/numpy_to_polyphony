module listc14r20_matmult (
    input wire clk,
    input wire rst,
    input wire matmult_ready,
    input wire matmult_accept,
    output reg matmult_valid,
    input wire signed [63:0] matmult_in_a0,
    input wire signed [63:0] matmult_in_a1,
    input wire signed [63:0] matmult_in_a2,
    input wire signed [63:0] matmult_in_a3,
    input wire signed [63:0] matmult_in_a4,
    input wire signed [63:0] matmult_in_a5,
    input wire signed [63:0] matmult_in_a6,
    input wire signed [63:0] matmult_in_a7,
    input wire signed [63:0] matmult_in_a8,
    input wire signed [63:0] matmult_in_a9,
    input wire signed [63:0] matmult_in_a10,
    input wire signed [63:0] matmult_in_a11,
    input wire signed [63:0] matmult_in_a12,
    input wire signed [63:0] matmult_in_a13,
    input wire signed [63:0] matmult_in_a14,
    input wire signed [63:0] matmult_in_a15,
    input wire signed [63:0] matmult_in_a16,
    input wire signed [63:0] matmult_in_a17,
    input wire signed [63:0] matmult_in_a18,
    input wire signed [63:0] matmult_in_a19,
    input wire signed [63:0] matmult_in_a20,
    input wire signed [63:0] matmult_in_a21,
    input wire signed [63:0] matmult_in_a22,
    input wire signed [63:0] matmult_in_a23,
    input wire signed [63:0] matmult_in_a24,
    input wire signed [63:0] matmult_in_a25,
    input wire signed [63:0] matmult_in_a26,
    input wire signed [63:0] matmult_in_a27,
    input wire signed [63:0] matmult_in_a28,
    input wire signed [63:0] matmult_in_a29,
    input wire signed [63:0] matmult_in_a30,
    input wire signed [63:0] matmult_in_a31,
    input wire signed [63:0] matmult_in_a32,
    input wire signed [63:0] matmult_in_a33,
    input wire signed [63:0] matmult_in_a34,
    input wire signed [63:0] matmult_in_a35,
    input wire signed [63:0] matmult_in_a36,
    input wire signed [63:0] matmult_in_a37,
    input wire signed [63:0] matmult_in_a38,
    input wire signed [63:0] matmult_in_a39,
    input wire signed [63:0] matmult_in_a40,
    input wire signed [63:0] matmult_in_a41,
    input wire signed [63:0] matmult_in_a42,
    input wire signed [63:0] matmult_in_a43,
    input wire signed [63:0] matmult_in_a44,
    input wire signed [63:0] matmult_in_a45,
    input wire signed [63:0] matmult_in_a46,
    input wire signed [63:0] matmult_in_a47,
    input wire signed [63:0] matmult_in_a48,
    input wire signed [63:0] matmult_in_a49,
    input wire signed [63:0] matmult_in_a50,
    input wire signed [63:0] matmult_in_a51,
    input wire signed [63:0] matmult_in_a52,
    input wire signed [63:0] matmult_in_a53,
    input wire signed [63:0] matmult_in_a54,
    input wire signed [63:0] matmult_in_a55,
    input wire signed [63:0] matmult_in_a56,
    input wire signed [63:0] matmult_in_a57,
    input wire signed [63:0] matmult_in_a58,
    input wire signed [63:0] matmult_in_a59,
    input wire signed [63:0] matmult_in_a60,
    input wire signed [63:0] matmult_in_a61,
    input wire signed [63:0] matmult_in_a62,
    input wire signed [63:0] matmult_in_a63,
    input wire signed [63:0] matmult_in_a64,
    input wire signed [63:0] matmult_in_a65,
    input wire signed [63:0] matmult_in_a66,
    input wire signed [63:0] matmult_in_a67,
    input wire signed [63:0] matmult_in_a68,
    input wire signed [63:0] matmult_in_a69,
    input wire signed [63:0] matmult_in_a70,
    input wire signed [63:0] matmult_in_a71,
    input wire signed [63:0] matmult_in_a72,
    input wire signed [63:0] matmult_in_a73,
    input wire signed [63:0] matmult_in_a74,
    input wire signed [63:0] matmult_in_a75,
    input wire signed [63:0] matmult_in_a76,
    input wire signed [63:0] matmult_in_a77,
    input wire signed [63:0] matmult_in_a78,
    input wire signed [63:0] matmult_in_a79,
    input wire signed [63:0] matmult_in_a80,
    input wire signed [63:0] matmult_in_a81,
    input wire signed [63:0] matmult_in_a82,
    input wire signed [63:0] matmult_in_a83,
    input wire signed [63:0] matmult_in_a84,
    input wire signed [63:0] matmult_in_a85,
    input wire signed [63:0] matmult_in_a86,
    input wire signed [63:0] matmult_in_a87,
    input wire signed [63:0] matmult_in_a88,
    input wire signed [63:0] matmult_in_a89,
    input wire signed [63:0] matmult_in_a90,
    input wire signed [63:0] matmult_in_a91,
    input wire signed [63:0] matmult_in_a92,
    input wire signed [63:0] matmult_in_a93,
    input wire signed [63:0] matmult_in_a94,
    input wire signed [63:0] matmult_in_a95,
    input wire signed [63:0] matmult_in_a96,
    input wire signed [63:0] matmult_in_a97,
    input wire signed [63:0] matmult_in_a98,
    input wire signed [63:0] matmult_in_a99,
    input wire signed [63:0] matmult_in_a100,
    input wire signed [63:0] matmult_in_a101,
    input wire signed [63:0] matmult_in_a102,
    input wire signed [63:0] matmult_in_a103,
    input wire signed [63:0] matmult_in_a104,
    input wire signed [63:0] matmult_in_a105,
    input wire signed [63:0] matmult_in_a106,
    input wire signed [63:0] matmult_in_a107,
    input wire signed [63:0] matmult_in_a108,
    input wire signed [63:0] matmult_in_a109,
    input wire signed [63:0] matmult_in_a110,
    input wire signed [63:0] matmult_in_a111,
    input wire signed [63:0] matmult_in_a112,
    input wire signed [63:0] matmult_in_a113,
    input wire signed [63:0] matmult_in_a114,
    input wire signed [63:0] matmult_in_a115,
    input wire signed [63:0] matmult_in_a116,
    input wire signed [63:0] matmult_in_a117,
    input wire signed [63:0] matmult_in_a118,
    input wire signed [63:0] matmult_in_a119,
    input wire signed [63:0] matmult_in_a120,
    input wire signed [63:0] matmult_in_a121,
    input wire signed [63:0] matmult_in_a122,
    input wire signed [63:0] matmult_in_a123,
    input wire signed [63:0] matmult_in_a124,
    input wire signed [63:0] matmult_in_a125,
    input wire signed [63:0] matmult_in_a126,
    input wire signed [63:0] matmult_in_a127,
    input wire signed [63:0] matmult_in_a128,
    input wire signed [63:0] matmult_in_a129,
    input wire signed [63:0] matmult_in_a130,
    input wire signed [63:0] matmult_in_a131,
    input wire signed [63:0] matmult_in_a132,
    input wire signed [63:0] matmult_in_a133,
    input wire signed [63:0] matmult_in_a134,
    input wire signed [63:0] matmult_in_a135,
    input wire signed [63:0] matmult_in_a136,
    input wire signed [63:0] matmult_in_a137,
    input wire signed [63:0] matmult_in_a138,
    input wire signed [63:0] matmult_in_a139,
    input wire signed [63:0] matmult_in_a140,
    input wire signed [63:0] matmult_in_a141,
    input wire signed [63:0] matmult_in_a142,
    input wire signed [63:0] matmult_in_a143,
    input wire signed [63:0] matmult_in_a144,
    input wire signed [63:0] matmult_in_a145,
    input wire signed [63:0] matmult_in_a146,
    input wire signed [63:0] matmult_in_a147,
    input wire signed [63:0] matmult_in_a148,
    input wire signed [63:0] matmult_in_a149,
    input wire signed [63:0] matmult_in_a150,
    input wire signed [63:0] matmult_in_a151,
    input wire signed [63:0] matmult_in_a152,
    input wire signed [63:0] matmult_in_a153,
    input wire signed [63:0] matmult_in_a154,
    input wire signed [63:0] matmult_in_a155,
    input wire signed [63:0] matmult_in_a156,
    input wire signed [63:0] matmult_in_a157,
    input wire signed [63:0] matmult_in_a158,
    input wire signed [63:0] matmult_in_a159,
    input wire signed [63:0] matmult_in_a160,
    input wire signed [63:0] matmult_in_a161,
    input wire signed [63:0] matmult_in_a162,
    input wire signed [63:0] matmult_in_a163,
    input wire signed [63:0] matmult_in_a164,
    input wire signed [63:0] matmult_in_a165,
    input wire signed [63:0] matmult_in_a166,
    input wire signed [63:0] matmult_in_a167,
    input wire signed [63:0] matmult_in_a168,
    input wire signed [63:0] matmult_in_a169,
    input wire signed [63:0] matmult_in_a170,
    input wire signed [63:0] matmult_in_a171,
    input wire signed [63:0] matmult_in_a172,
    input wire signed [63:0] matmult_in_a173,
    input wire signed [63:0] matmult_in_a174,
    input wire signed [63:0] matmult_in_a175,
    input wire signed [63:0] matmult_in_a176,
    input wire signed [63:0] matmult_in_a177,
    input wire signed [63:0] matmult_in_a178,
    input wire signed [63:0] matmult_in_a179,
    input wire signed [63:0] matmult_in_a180,
    input wire signed [63:0] matmult_in_a181,
    input wire signed [63:0] matmult_in_a182,
    input wire signed [63:0] matmult_in_a183,
    input wire signed [63:0] matmult_in_a184,
    input wire signed [63:0] matmult_in_a185,
    input wire signed [63:0] matmult_in_a186,
    input wire signed [63:0] matmult_in_a187,
    input wire signed [63:0] matmult_in_a188,
    input wire signed [63:0] matmult_in_a189,
    input wire signed [63:0] matmult_in_a190,
    input wire signed [63:0] matmult_in_a191,
    input wire signed [63:0] matmult_in_a192,
    input wire signed [63:0] matmult_in_a193,
    input wire signed [63:0] matmult_in_a194,
    input wire signed [63:0] matmult_in_a195,
    input wire signed [63:0] matmult_in_a196,
    input wire signed [63:0] matmult_in_a197,
    input wire signed [63:0] matmult_in_a198,
    input wire signed [63:0] matmult_in_a199,
    input wire signed [63:0] matmult_in_a200,
    input wire signed [63:0] matmult_in_a201,
    input wire signed [63:0] matmult_in_a202,
    input wire signed [63:0] matmult_in_a203,
    input wire signed [63:0] matmult_in_a204,
    input wire signed [63:0] matmult_in_a205,
    input wire signed [63:0] matmult_in_a206,
    input wire signed [63:0] matmult_in_a207,
    input wire signed [63:0] matmult_in_a208,
    input wire signed [63:0] matmult_in_a209,
    input wire signed [63:0] matmult_in_a210,
    input wire signed [63:0] matmult_in_a211,
    input wire signed [63:0] matmult_in_a212,
    input wire signed [63:0] matmult_in_a213,
    input wire signed [63:0] matmult_in_a214,
    input wire signed [63:0] matmult_in_a215,
    input wire signed [63:0] matmult_in_a216,
    input wire signed [63:0] matmult_in_a217,
    input wire signed [63:0] matmult_in_a218,
    input wire signed [63:0] matmult_in_a219,
    input wire signed [63:0] matmult_in_a220,
    input wire signed [63:0] matmult_in_a221,
    input wire signed [63:0] matmult_in_a222,
    input wire signed [63:0] matmult_in_a223,
    input wire signed [63:0] matmult_in_a224,
    input wire signed [63:0] matmult_in_a225,
    input wire signed [63:0] matmult_in_a226,
    input wire signed [63:0] matmult_in_a227,
    input wire signed [63:0] matmult_in_a228,
    input wire signed [63:0] matmult_in_a229,
    input wire signed [63:0] matmult_in_a230,
    input wire signed [63:0] matmult_in_a231,
    input wire signed [63:0] matmult_in_a232,
    input wire signed [63:0] matmult_in_a233,
    input wire signed [63:0] matmult_in_a234,
    input wire signed [63:0] matmult_in_a235,
    input wire signed [63:0] matmult_in_a236,
    input wire signed [63:0] matmult_in_a237,
    input wire signed [63:0] matmult_in_a238,
    input wire signed [63:0] matmult_in_a239,
    input wire signed [63:0] matmult_in_a240,
    input wire signed [63:0] matmult_in_a241,
    input wire signed [63:0] matmult_in_a242,
    input wire signed [63:0] matmult_in_a243,
    input wire signed [63:0] matmult_in_a244,
    input wire signed [63:0] matmult_in_a245,
    input wire signed [63:0] matmult_in_a246,
    input wire signed [63:0] matmult_in_a247,
    input wire signed [63:0] matmult_in_a248,
    input wire signed [63:0] matmult_in_a249,
    input wire signed [63:0] matmult_in_a250,
    input wire signed [63:0] matmult_in_a251,
    input wire signed [63:0] matmult_in_a252,
    input wire signed [63:0] matmult_in_a253,
    input wire signed [63:0] matmult_in_a254,
    input wire signed [63:0] matmult_in_a255,
    input wire signed [63:0] matmult_in_a256,
    input wire signed [63:0] matmult_in_a257,
    input wire signed [63:0] matmult_in_a258,
    input wire signed [63:0] matmult_in_a259,
    input wire signed [63:0] matmult_in_a260,
    input wire signed [63:0] matmult_in_a261,
    input wire signed [63:0] matmult_in_a262,
    input wire signed [63:0] matmult_in_a263,
    input wire signed [63:0] matmult_in_a264,
    input wire signed [63:0] matmult_in_a265,
    input wire signed [63:0] matmult_in_a266,
    input wire signed [63:0] matmult_in_a267,
    input wire signed [63:0] matmult_in_a268,
    input wire signed [63:0] matmult_in_a269,
    input wire signed [63:0] matmult_in_a270,
    input wire signed [63:0] matmult_in_a271,
    input wire signed [63:0] matmult_in_a272,
    input wire signed [63:0] matmult_in_a273,
    input wire signed [63:0] matmult_in_a274,
    input wire signed [63:0] matmult_in_a275,
    input wire signed [63:0] matmult_in_a276,
    input wire signed [63:0] matmult_in_a277,
    input wire signed [63:0] matmult_in_a278,
    input wire signed [63:0] matmult_in_a279,
    output wire signed [63:0] matmult_out_a0,
    output wire signed [63:0] matmult_out_a1,
    output wire signed [63:0] matmult_out_a2,
    output wire signed [63:0] matmult_out_a3,
    output wire signed [63:0] matmult_out_a4,
    output wire signed [63:0] matmult_out_a5,
    output wire signed [63:0] matmult_out_a6,
    output wire signed [63:0] matmult_out_a7,
    output wire signed [63:0] matmult_out_a8,
    output wire signed [63:0] matmult_out_a9,
    output wire signed [63:0] matmult_out_a10,
    output wire signed [63:0] matmult_out_a11,
    output wire signed [63:0] matmult_out_a12,
    output wire signed [63:0] matmult_out_a13,
    output wire signed [63:0] matmult_out_a14,
    output wire signed [63:0] matmult_out_a15,
    output wire signed [63:0] matmult_out_a16,
    output wire signed [63:0] matmult_out_a17,
    output wire signed [63:0] matmult_out_a18,
    output wire signed [63:0] matmult_out_a19,
    output wire signed [63:0] matmult_out_a20,
    output wire signed [63:0] matmult_out_a21,
    output wire signed [63:0] matmult_out_a22,
    output wire signed [63:0] matmult_out_a23,
    output wire signed [63:0] matmult_out_a24,
    output wire signed [63:0] matmult_out_a25,
    output wire signed [63:0] matmult_out_a26,
    output wire signed [63:0] matmult_out_a27,
    output wire signed [63:0] matmult_out_a28,
    output wire signed [63:0] matmult_out_a29,
    output wire signed [63:0] matmult_out_a30,
    output wire signed [63:0] matmult_out_a31,
    output wire signed [63:0] matmult_out_a32,
    output wire signed [63:0] matmult_out_a33,
    output wire signed [63:0] matmult_out_a34,
    output wire signed [63:0] matmult_out_a35,
    output wire signed [63:0] matmult_out_a36,
    output wire signed [63:0] matmult_out_a37,
    output wire signed [63:0] matmult_out_a38,
    output wire signed [63:0] matmult_out_a39,
    output wire signed [63:0] matmult_out_a40,
    output wire signed [63:0] matmult_out_a41,
    output wire signed [63:0] matmult_out_a42,
    output wire signed [63:0] matmult_out_a43,
    output wire signed [63:0] matmult_out_a44,
    output wire signed [63:0] matmult_out_a45,
    output wire signed [63:0] matmult_out_a46,
    output wire signed [63:0] matmult_out_a47,
    output wire signed [63:0] matmult_out_a48,
    output wire signed [63:0] matmult_out_a49,
    output wire signed [63:0] matmult_out_a50,
    output wire signed [63:0] matmult_out_a51,
    output wire signed [63:0] matmult_out_a52,
    output wire signed [63:0] matmult_out_a53,
    output wire signed [63:0] matmult_out_a54,
    output wire signed [63:0] matmult_out_a55,
    output wire signed [63:0] matmult_out_a56,
    output wire signed [63:0] matmult_out_a57,
    output wire signed [63:0] matmult_out_a58,
    output wire signed [63:0] matmult_out_a59,
    output wire signed [63:0] matmult_out_a60,
    output wire signed [63:0] matmult_out_a61,
    output wire signed [63:0] matmult_out_a62,
    output wire signed [63:0] matmult_out_a63,
    output wire signed [63:0] matmult_out_a64,
    output wire signed [63:0] matmult_out_a65,
    output wire signed [63:0] matmult_out_a66,
    output wire signed [63:0] matmult_out_a67,
    output wire signed [63:0] matmult_out_a68,
    output wire signed [63:0] matmult_out_a69,
    output wire signed [63:0] matmult_out_a70,
    output wire signed [63:0] matmult_out_a71,
    output wire signed [63:0] matmult_out_a72,
    output wire signed [63:0] matmult_out_a73,
    output wire signed [63:0] matmult_out_a74,
    output wire signed [63:0] matmult_out_a75,
    output wire signed [63:0] matmult_out_a76,
    output wire signed [63:0] matmult_out_a77,
    output wire signed [63:0] matmult_out_a78,
    output wire signed [63:0] matmult_out_a79,
    output wire signed [63:0] matmult_out_a80,
    output wire signed [63:0] matmult_out_a81,
    output wire signed [63:0] matmult_out_a82,
    output wire signed [63:0] matmult_out_a83,
    output wire signed [63:0] matmult_out_a84,
    output wire signed [63:0] matmult_out_a85,
    output wire signed [63:0] matmult_out_a86,
    output wire signed [63:0] matmult_out_a87,
    output wire signed [63:0] matmult_out_a88,
    output wire signed [63:0] matmult_out_a89,
    output wire signed [63:0] matmult_out_a90,
    output wire signed [63:0] matmult_out_a91,
    output wire signed [63:0] matmult_out_a92,
    output wire signed [63:0] matmult_out_a93,
    output wire signed [63:0] matmult_out_a94,
    output wire signed [63:0] matmult_out_a95,
    output wire signed [63:0] matmult_out_a96,
    output wire signed [63:0] matmult_out_a97,
    output wire signed [63:0] matmult_out_a98,
    output wire signed [63:0] matmult_out_a99,
    output wire signed [63:0] matmult_out_a100,
    output wire signed [63:0] matmult_out_a101,
    output wire signed [63:0] matmult_out_a102,
    output wire signed [63:0] matmult_out_a103,
    output wire signed [63:0] matmult_out_a104,
    output wire signed [63:0] matmult_out_a105,
    output wire signed [63:0] matmult_out_a106,
    output wire signed [63:0] matmult_out_a107,
    output wire signed [63:0] matmult_out_a108,
    output wire signed [63:0] matmult_out_a109,
    output wire signed [63:0] matmult_out_a110,
    output wire signed [63:0] matmult_out_a111,
    output wire signed [63:0] matmult_out_a112,
    output wire signed [63:0] matmult_out_a113,
    output wire signed [63:0] matmult_out_a114,
    output wire signed [63:0] matmult_out_a115,
    output wire signed [63:0] matmult_out_a116,
    output wire signed [63:0] matmult_out_a117,
    output wire signed [63:0] matmult_out_a118,
    output wire signed [63:0] matmult_out_a119,
    output wire signed [63:0] matmult_out_a120,
    output wire signed [63:0] matmult_out_a121,
    output wire signed [63:0] matmult_out_a122,
    output wire signed [63:0] matmult_out_a123,
    output wire signed [63:0] matmult_out_a124,
    output wire signed [63:0] matmult_out_a125,
    output wire signed [63:0] matmult_out_a126,
    output wire signed [63:0] matmult_out_a127,
    output wire signed [63:0] matmult_out_a128,
    output wire signed [63:0] matmult_out_a129,
    output wire signed [63:0] matmult_out_a130,
    output wire signed [63:0] matmult_out_a131,
    output wire signed [63:0] matmult_out_a132,
    output wire signed [63:0] matmult_out_a133,
    output wire signed [63:0] matmult_out_a134,
    output wire signed [63:0] matmult_out_a135,
    output wire signed [63:0] matmult_out_a136,
    output wire signed [63:0] matmult_out_a137,
    output wire signed [63:0] matmult_out_a138,
    output wire signed [63:0] matmult_out_a139,
    output wire signed [63:0] matmult_out_a140,
    output wire signed [63:0] matmult_out_a141,
    output wire signed [63:0] matmult_out_a142,
    output wire signed [63:0] matmult_out_a143,
    output wire signed [63:0] matmult_out_a144,
    output wire signed [63:0] matmult_out_a145,
    output wire signed [63:0] matmult_out_a146,
    output wire signed [63:0] matmult_out_a147,
    output wire signed [63:0] matmult_out_a148,
    output wire signed [63:0] matmult_out_a149,
    output wire signed [63:0] matmult_out_a150,
    output wire signed [63:0] matmult_out_a151,
    output wire signed [63:0] matmult_out_a152,
    output wire signed [63:0] matmult_out_a153,
    output wire signed [63:0] matmult_out_a154,
    output wire signed [63:0] matmult_out_a155,
    output wire signed [63:0] matmult_out_a156,
    output wire signed [63:0] matmult_out_a157,
    output wire signed [63:0] matmult_out_a158,
    output wire signed [63:0] matmult_out_a159,
    output wire signed [63:0] matmult_out_a160,
    output wire signed [63:0] matmult_out_a161,
    output wire signed [63:0] matmult_out_a162,
    output wire signed [63:0] matmult_out_a163,
    output wire signed [63:0] matmult_out_a164,
    output wire signed [63:0] matmult_out_a165,
    output wire signed [63:0] matmult_out_a166,
    output wire signed [63:0] matmult_out_a167,
    output wire signed [63:0] matmult_out_a168,
    output wire signed [63:0] matmult_out_a169,
    output wire signed [63:0] matmult_out_a170,
    output wire signed [63:0] matmult_out_a171,
    output wire signed [63:0] matmult_out_a172,
    output wire signed [63:0] matmult_out_a173,
    output wire signed [63:0] matmult_out_a174,
    output wire signed [63:0] matmult_out_a175,
    output wire signed [63:0] matmult_out_a176,
    output wire signed [63:0] matmult_out_a177,
    output wire signed [63:0] matmult_out_a178,
    output wire signed [63:0] matmult_out_a179,
    output wire signed [63:0] matmult_out_a180,
    output wire signed [63:0] matmult_out_a181,
    output wire signed [63:0] matmult_out_a182,
    output wire signed [63:0] matmult_out_a183,
    output wire signed [63:0] matmult_out_a184,
    output wire signed [63:0] matmult_out_a185,
    output wire signed [63:0] matmult_out_a186,
    output wire signed [63:0] matmult_out_a187,
    output wire signed [63:0] matmult_out_a188,
    output wire signed [63:0] matmult_out_a189,
    output wire signed [63:0] matmult_out_a190,
    output wire signed [63:0] matmult_out_a191,
    output wire signed [63:0] matmult_out_a192,
    output wire signed [63:0] matmult_out_a193,
    output wire signed [63:0] matmult_out_a194,
    output wire signed [63:0] matmult_out_a195,
    output wire signed [63:0] matmult_out_a196,
    output wire signed [63:0] matmult_out_a197,
    output wire signed [63:0] matmult_out_a198,
    output wire signed [63:0] matmult_out_a199,
    output wire signed [63:0] matmult_out_a200,
    output wire signed [63:0] matmult_out_a201,
    output wire signed [63:0] matmult_out_a202,
    output wire signed [63:0] matmult_out_a203,
    output wire signed [63:0] matmult_out_a204,
    output wire signed [63:0] matmult_out_a205,
    output wire signed [63:0] matmult_out_a206,
    output wire signed [63:0] matmult_out_a207,
    output wire signed [63:0] matmult_out_a208,
    output wire signed [63:0] matmult_out_a209,
    output wire signed [63:0] matmult_out_a210,
    output wire signed [63:0] matmult_out_a211,
    output wire signed [63:0] matmult_out_a212,
    output wire signed [63:0] matmult_out_a213,
    output wire signed [63:0] matmult_out_a214,
    output wire signed [63:0] matmult_out_a215,
    output wire signed [63:0] matmult_out_a216,
    output wire signed [63:0] matmult_out_a217,
    output wire signed [63:0] matmult_out_a218,
    output wire signed [63:0] matmult_out_a219,
    output wire signed [63:0] matmult_out_a220,
    output wire signed [63:0] matmult_out_a221,
    output wire signed [63:0] matmult_out_a222,
    output wire signed [63:0] matmult_out_a223,
    output wire signed [63:0] matmult_out_a224,
    output wire signed [63:0] matmult_out_a225,
    output wire signed [63:0] matmult_out_a226,
    output wire signed [63:0] matmult_out_a227,
    output wire signed [63:0] matmult_out_a228,
    output wire signed [63:0] matmult_out_a229,
    output wire signed [63:0] matmult_out_a230,
    output wire signed [63:0] matmult_out_a231,
    output wire signed [63:0] matmult_out_a232,
    output wire signed [63:0] matmult_out_a233,
    output wire signed [63:0] matmult_out_a234,
    output wire signed [63:0] matmult_out_a235,
    output wire signed [63:0] matmult_out_a236,
    output wire signed [63:0] matmult_out_a237,
    output wire signed [63:0] matmult_out_a238,
    output wire signed [63:0] matmult_out_a239,
    output wire signed [63:0] matmult_out_a240,
    output wire signed [63:0] matmult_out_a241,
    output wire signed [63:0] matmult_out_a242,
    output wire signed [63:0] matmult_out_a243,
    output wire signed [63:0] matmult_out_a244,
    output wire signed [63:0] matmult_out_a245,
    output wire signed [63:0] matmult_out_a246,
    output wire signed [63:0] matmult_out_a247,
    output wire signed [63:0] matmult_out_a248,
    output wire signed [63:0] matmult_out_a249,
    output wire signed [63:0] matmult_out_a250,
    output wire signed [63:0] matmult_out_a251,
    output wire signed [63:0] matmult_out_a252,
    output wire signed [63:0] matmult_out_a253,
    output wire signed [63:0] matmult_out_a254,
    output wire signed [63:0] matmult_out_a255,
    output wire signed [63:0] matmult_out_a256,
    output wire signed [63:0] matmult_out_a257,
    output wire signed [63:0] matmult_out_a258,
    output wire signed [63:0] matmult_out_a259,
    output wire signed [63:0] matmult_out_a260,
    output wire signed [63:0] matmult_out_a261,
    output wire signed [63:0] matmult_out_a262,
    output wire signed [63:0] matmult_out_a263,
    output wire signed [63:0] matmult_out_a264,
    output wire signed [63:0] matmult_out_a265,
    output wire signed [63:0] matmult_out_a266,
    output wire signed [63:0] matmult_out_a267,
    output wire signed [63:0] matmult_out_a268,
    output wire signed [63:0] matmult_out_a269,
    output wire signed [63:0] matmult_out_a270,
    output wire signed [63:0] matmult_out_a271,
    output wire signed [63:0] matmult_out_a272,
    output wire signed [63:0] matmult_out_a273,
    output wire signed [63:0] matmult_out_a274,
    output wire signed [63:0] matmult_out_a275,
    output wire signed [63:0] matmult_out_a276,
    output wire signed [63:0] matmult_out_a277,
    output wire signed [63:0] matmult_out_a278,
    output wire signed [63:0] matmult_out_a279,
    input wire signed [63:0] matmult_in_b0,
    input wire signed [63:0] matmult_in_b1,
    input wire signed [63:0] matmult_in_b2,
    input wire signed [63:0] matmult_in_b3,
    input wire signed [63:0] matmult_in_b4,
    input wire signed [63:0] matmult_in_b5,
    input wire signed [63:0] matmult_in_b6,
    input wire signed [63:0] matmult_in_b7,
    input wire signed [63:0] matmult_in_b8,
    input wire signed [63:0] matmult_in_b9,
    input wire signed [63:0] matmult_in_b10,
    input wire signed [63:0] matmult_in_b11,
    input wire signed [63:0] matmult_in_b12,
    input wire signed [63:0] matmult_in_b13,
    input wire signed [63:0] matmult_in_b14,
    input wire signed [63:0] matmult_in_b15,
    input wire signed [63:0] matmult_in_b16,
    input wire signed [63:0] matmult_in_b17,
    input wire signed [63:0] matmult_in_b18,
    input wire signed [63:0] matmult_in_b19,
    input wire signed [63:0] matmult_in_b20,
    input wire signed [63:0] matmult_in_b21,
    input wire signed [63:0] matmult_in_b22,
    input wire signed [63:0] matmult_in_b23,
    input wire signed [63:0] matmult_in_b24,
    input wire signed [63:0] matmult_in_b25,
    input wire signed [63:0] matmult_in_b26,
    input wire signed [63:0] matmult_in_b27,
    input wire signed [63:0] matmult_in_b28,
    input wire signed [63:0] matmult_in_b29,
    input wire signed [63:0] matmult_in_b30,
    input wire signed [63:0] matmult_in_b31,
    input wire signed [63:0] matmult_in_b32,
    input wire signed [63:0] matmult_in_b33,
    input wire signed [63:0] matmult_in_b34,
    input wire signed [63:0] matmult_in_b35,
    input wire signed [63:0] matmult_in_b36,
    input wire signed [63:0] matmult_in_b37,
    input wire signed [63:0] matmult_in_b38,
    input wire signed [63:0] matmult_in_b39,
    input wire signed [63:0] matmult_in_b40,
    input wire signed [63:0] matmult_in_b41,
    input wire signed [63:0] matmult_in_b42,
    input wire signed [63:0] matmult_in_b43,
    input wire signed [63:0] matmult_in_b44,
    input wire signed [63:0] matmult_in_b45,
    input wire signed [63:0] matmult_in_b46,
    input wire signed [63:0] matmult_in_b47,
    input wire signed [63:0] matmult_in_b48,
    input wire signed [63:0] matmult_in_b49,
    input wire signed [63:0] matmult_in_b50,
    input wire signed [63:0] matmult_in_b51,
    input wire signed [63:0] matmult_in_b52,
    input wire signed [63:0] matmult_in_b53,
    input wire signed [63:0] matmult_in_b54,
    input wire signed [63:0] matmult_in_b55,
    input wire signed [63:0] matmult_in_b56,
    input wire signed [63:0] matmult_in_b57,
    input wire signed [63:0] matmult_in_b58,
    input wire signed [63:0] matmult_in_b59,
    input wire signed [63:0] matmult_in_b60,
    input wire signed [63:0] matmult_in_b61,
    input wire signed [63:0] matmult_in_b62,
    input wire signed [63:0] matmult_in_b63,
    input wire signed [63:0] matmult_in_b64,
    input wire signed [63:0] matmult_in_b65,
    input wire signed [63:0] matmult_in_b66,
    input wire signed [63:0] matmult_in_b67,
    input wire signed [63:0] matmult_in_b68,
    input wire signed [63:0] matmult_in_b69,
    input wire signed [63:0] matmult_in_b70,
    input wire signed [63:0] matmult_in_b71,
    input wire signed [63:0] matmult_in_b72,
    input wire signed [63:0] matmult_in_b73,
    input wire signed [63:0] matmult_in_b74,
    input wire signed [63:0] matmult_in_b75,
    input wire signed [63:0] matmult_in_b76,
    input wire signed [63:0] matmult_in_b77,
    input wire signed [63:0] matmult_in_b78,
    input wire signed [63:0] matmult_in_b79,
    input wire signed [63:0] matmult_in_b80,
    input wire signed [63:0] matmult_in_b81,
    input wire signed [63:0] matmult_in_b82,
    input wire signed [63:0] matmult_in_b83,
    input wire signed [63:0] matmult_in_b84,
    input wire signed [63:0] matmult_in_b85,
    input wire signed [63:0] matmult_in_b86,
    input wire signed [63:0] matmult_in_b87,
    input wire signed [63:0] matmult_in_b88,
    input wire signed [63:0] matmult_in_b89,
    input wire signed [63:0] matmult_in_b90,
    input wire signed [63:0] matmult_in_b91,
    input wire signed [63:0] matmult_in_b92,
    input wire signed [63:0] matmult_in_b93,
    input wire signed [63:0] matmult_in_b94,
    input wire signed [63:0] matmult_in_b95,
    input wire signed [63:0] matmult_in_b96,
    input wire signed [63:0] matmult_in_b97,
    input wire signed [63:0] matmult_in_b98,
    input wire signed [63:0] matmult_in_b99,
    input wire signed [63:0] matmult_in_b100,
    input wire signed [63:0] matmult_in_b101,
    input wire signed [63:0] matmult_in_b102,
    input wire signed [63:0] matmult_in_b103,
    input wire signed [63:0] matmult_in_b104,
    input wire signed [63:0] matmult_in_b105,
    input wire signed [63:0] matmult_in_b106,
    input wire signed [63:0] matmult_in_b107,
    input wire signed [63:0] matmult_in_b108,
    input wire signed [63:0] matmult_in_b109,
    input wire signed [63:0] matmult_in_b110,
    input wire signed [63:0] matmult_in_b111,
    input wire signed [63:0] matmult_in_b112,
    input wire signed [63:0] matmult_in_b113,
    input wire signed [63:0] matmult_in_b114,
    input wire signed [63:0] matmult_in_b115,
    input wire signed [63:0] matmult_in_b116,
    input wire signed [63:0] matmult_in_b117,
    input wire signed [63:0] matmult_in_b118,
    input wire signed [63:0] matmult_in_b119,
    input wire signed [63:0] matmult_in_b120,
    input wire signed [63:0] matmult_in_b121,
    input wire signed [63:0] matmult_in_b122,
    input wire signed [63:0] matmult_in_b123,
    input wire signed [63:0] matmult_in_b124,
    input wire signed [63:0] matmult_in_b125,
    input wire signed [63:0] matmult_in_b126,
    input wire signed [63:0] matmult_in_b127,
    input wire signed [63:0] matmult_in_b128,
    input wire signed [63:0] matmult_in_b129,
    input wire signed [63:0] matmult_in_b130,
    input wire signed [63:0] matmult_in_b131,
    input wire signed [63:0] matmult_in_b132,
    input wire signed [63:0] matmult_in_b133,
    input wire signed [63:0] matmult_in_b134,
    input wire signed [63:0] matmult_in_b135,
    input wire signed [63:0] matmult_in_b136,
    input wire signed [63:0] matmult_in_b137,
    input wire signed [63:0] matmult_in_b138,
    input wire signed [63:0] matmult_in_b139,
    input wire signed [63:0] matmult_in_b140,
    input wire signed [63:0] matmult_in_b141,
    input wire signed [63:0] matmult_in_b142,
    input wire signed [63:0] matmult_in_b143,
    input wire signed [63:0] matmult_in_b144,
    input wire signed [63:0] matmult_in_b145,
    input wire signed [63:0] matmult_in_b146,
    input wire signed [63:0] matmult_in_b147,
    input wire signed [63:0] matmult_in_b148,
    input wire signed [63:0] matmult_in_b149,
    input wire signed [63:0] matmult_in_b150,
    input wire signed [63:0] matmult_in_b151,
    input wire signed [63:0] matmult_in_b152,
    input wire signed [63:0] matmult_in_b153,
    input wire signed [63:0] matmult_in_b154,
    input wire signed [63:0] matmult_in_b155,
    input wire signed [63:0] matmult_in_b156,
    input wire signed [63:0] matmult_in_b157,
    input wire signed [63:0] matmult_in_b158,
    input wire signed [63:0] matmult_in_b159,
    input wire signed [63:0] matmult_in_b160,
    input wire signed [63:0] matmult_in_b161,
    input wire signed [63:0] matmult_in_b162,
    input wire signed [63:0] matmult_in_b163,
    input wire signed [63:0] matmult_in_b164,
    input wire signed [63:0] matmult_in_b165,
    input wire signed [63:0] matmult_in_b166,
    input wire signed [63:0] matmult_in_b167,
    input wire signed [63:0] matmult_in_b168,
    input wire signed [63:0] matmult_in_b169,
    input wire signed [63:0] matmult_in_b170,
    input wire signed [63:0] matmult_in_b171,
    input wire signed [63:0] matmult_in_b172,
    input wire signed [63:0] matmult_in_b173,
    input wire signed [63:0] matmult_in_b174,
    input wire signed [63:0] matmult_in_b175,
    input wire signed [63:0] matmult_in_b176,
    input wire signed [63:0] matmult_in_b177,
    input wire signed [63:0] matmult_in_b178,
    input wire signed [63:0] matmult_in_b179,
    input wire signed [63:0] matmult_in_b180,
    input wire signed [63:0] matmult_in_b181,
    input wire signed [63:0] matmult_in_b182,
    input wire signed [63:0] matmult_in_b183,
    input wire signed [63:0] matmult_in_b184,
    input wire signed [63:0] matmult_in_b185,
    input wire signed [63:0] matmult_in_b186,
    input wire signed [63:0] matmult_in_b187,
    input wire signed [63:0] matmult_in_b188,
    input wire signed [63:0] matmult_in_b189,
    input wire signed [63:0] matmult_in_b190,
    input wire signed [63:0] matmult_in_b191,
    input wire signed [63:0] matmult_in_b192,
    input wire signed [63:0] matmult_in_b193,
    input wire signed [63:0] matmult_in_b194,
    input wire signed [63:0] matmult_in_b195,
    input wire signed [63:0] matmult_in_b196,
    input wire signed [63:0] matmult_in_b197,
    input wire signed [63:0] matmult_in_b198,
    input wire signed [63:0] matmult_in_b199,
    input wire signed [63:0] matmult_in_b200,
    input wire signed [63:0] matmult_in_b201,
    input wire signed [63:0] matmult_in_b202,
    input wire signed [63:0] matmult_in_b203,
    input wire signed [63:0] matmult_in_b204,
    input wire signed [63:0] matmult_in_b205,
    input wire signed [63:0] matmult_in_b206,
    input wire signed [63:0] matmult_in_b207,
    input wire signed [63:0] matmult_in_b208,
    input wire signed [63:0] matmult_in_b209,
    input wire signed [63:0] matmult_in_b210,
    input wire signed [63:0] matmult_in_b211,
    input wire signed [63:0] matmult_in_b212,
    input wire signed [63:0] matmult_in_b213,
    input wire signed [63:0] matmult_in_b214,
    input wire signed [63:0] matmult_in_b215,
    input wire signed [63:0] matmult_in_b216,
    input wire signed [63:0] matmult_in_b217,
    input wire signed [63:0] matmult_in_b218,
    input wire signed [63:0] matmult_in_b219,
    input wire signed [63:0] matmult_in_b220,
    input wire signed [63:0] matmult_in_b221,
    input wire signed [63:0] matmult_in_b222,
    input wire signed [63:0] matmult_in_b223,
    input wire signed [63:0] matmult_in_b224,
    input wire signed [63:0] matmult_in_b225,
    input wire signed [63:0] matmult_in_b226,
    input wire signed [63:0] matmult_in_b227,
    input wire signed [63:0] matmult_in_b228,
    input wire signed [63:0] matmult_in_b229,
    input wire signed [63:0] matmult_in_b230,
    input wire signed [63:0] matmult_in_b231,
    input wire signed [63:0] matmult_in_b232,
    input wire signed [63:0] matmult_in_b233,
    input wire signed [63:0] matmult_in_b234,
    input wire signed [63:0] matmult_in_b235,
    input wire signed [63:0] matmult_in_b236,
    input wire signed [63:0] matmult_in_b237,
    input wire signed [63:0] matmult_in_b238,
    input wire signed [63:0] matmult_in_b239,
    input wire signed [63:0] matmult_in_b240,
    input wire signed [63:0] matmult_in_b241,
    input wire signed [63:0] matmult_in_b242,
    input wire signed [63:0] matmult_in_b243,
    input wire signed [63:0] matmult_in_b244,
    input wire signed [63:0] matmult_in_b245,
    input wire signed [63:0] matmult_in_b246,
    input wire signed [63:0] matmult_in_b247,
    input wire signed [63:0] matmult_in_b248,
    input wire signed [63:0] matmult_in_b249,
    input wire signed [63:0] matmult_in_b250,
    input wire signed [63:0] matmult_in_b251,
    input wire signed [63:0] matmult_in_b252,
    input wire signed [63:0] matmult_in_b253,
    input wire signed [63:0] matmult_in_b254,
    input wire signed [63:0] matmult_in_b255,
    input wire signed [63:0] matmult_in_b256,
    input wire signed [63:0] matmult_in_b257,
    input wire signed [63:0] matmult_in_b258,
    input wire signed [63:0] matmult_in_b259,
    input wire signed [63:0] matmult_in_b260,
    input wire signed [63:0] matmult_in_b261,
    input wire signed [63:0] matmult_in_b262,
    input wire signed [63:0] matmult_in_b263,
    input wire signed [63:0] matmult_in_b264,
    input wire signed [63:0] matmult_in_b265,
    input wire signed [63:0] matmult_in_b266,
    input wire signed [63:0] matmult_in_b267,
    input wire signed [63:0] matmult_in_b268,
    input wire signed [63:0] matmult_in_b269,
    input wire signed [63:0] matmult_in_b270,
    input wire signed [63:0] matmult_in_b271,
    input wire signed [63:0] matmult_in_b272,
    input wire signed [63:0] matmult_in_b273,
    input wire signed [63:0] matmult_in_b274,
    input wire signed [63:0] matmult_in_b275,
    input wire signed [63:0] matmult_in_b276,
    input wire signed [63:0] matmult_in_b277,
    input wire signed [63:0] matmult_in_b278,
    input wire signed [63:0] matmult_in_b279,
    output wire signed [63:0] matmult_out_b0,
    output wire signed [63:0] matmult_out_b1,
    output wire signed [63:0] matmult_out_b2,
    output wire signed [63:0] matmult_out_b3,
    output wire signed [63:0] matmult_out_b4,
    output wire signed [63:0] matmult_out_b5,
    output wire signed [63:0] matmult_out_b6,
    output wire signed [63:0] matmult_out_b7,
    output wire signed [63:0] matmult_out_b8,
    output wire signed [63:0] matmult_out_b9,
    output wire signed [63:0] matmult_out_b10,
    output wire signed [63:0] matmult_out_b11,
    output wire signed [63:0] matmult_out_b12,
    output wire signed [63:0] matmult_out_b13,
    output wire signed [63:0] matmult_out_b14,
    output wire signed [63:0] matmult_out_b15,
    output wire signed [63:0] matmult_out_b16,
    output wire signed [63:0] matmult_out_b17,
    output wire signed [63:0] matmult_out_b18,
    output wire signed [63:0] matmult_out_b19,
    output wire signed [63:0] matmult_out_b20,
    output wire signed [63:0] matmult_out_b21,
    output wire signed [63:0] matmult_out_b22,
    output wire signed [63:0] matmult_out_b23,
    output wire signed [63:0] matmult_out_b24,
    output wire signed [63:0] matmult_out_b25,
    output wire signed [63:0] matmult_out_b26,
    output wire signed [63:0] matmult_out_b27,
    output wire signed [63:0] matmult_out_b28,
    output wire signed [63:0] matmult_out_b29,
    output wire signed [63:0] matmult_out_b30,
    output wire signed [63:0] matmult_out_b31,
    output wire signed [63:0] matmult_out_b32,
    output wire signed [63:0] matmult_out_b33,
    output wire signed [63:0] matmult_out_b34,
    output wire signed [63:0] matmult_out_b35,
    output wire signed [63:0] matmult_out_b36,
    output wire signed [63:0] matmult_out_b37,
    output wire signed [63:0] matmult_out_b38,
    output wire signed [63:0] matmult_out_b39,
    output wire signed [63:0] matmult_out_b40,
    output wire signed [63:0] matmult_out_b41,
    output wire signed [63:0] matmult_out_b42,
    output wire signed [63:0] matmult_out_b43,
    output wire signed [63:0] matmult_out_b44,
    output wire signed [63:0] matmult_out_b45,
    output wire signed [63:0] matmult_out_b46,
    output wire signed [63:0] matmult_out_b47,
    output wire signed [63:0] matmult_out_b48,
    output wire signed [63:0] matmult_out_b49,
    output wire signed [63:0] matmult_out_b50,
    output wire signed [63:0] matmult_out_b51,
    output wire signed [63:0] matmult_out_b52,
    output wire signed [63:0] matmult_out_b53,
    output wire signed [63:0] matmult_out_b54,
    output wire signed [63:0] matmult_out_b55,
    output wire signed [63:0] matmult_out_b56,
    output wire signed [63:0] matmult_out_b57,
    output wire signed [63:0] matmult_out_b58,
    output wire signed [63:0] matmult_out_b59,
    output wire signed [63:0] matmult_out_b60,
    output wire signed [63:0] matmult_out_b61,
    output wire signed [63:0] matmult_out_b62,
    output wire signed [63:0] matmult_out_b63,
    output wire signed [63:0] matmult_out_b64,
    output wire signed [63:0] matmult_out_b65,
    output wire signed [63:0] matmult_out_b66,
    output wire signed [63:0] matmult_out_b67,
    output wire signed [63:0] matmult_out_b68,
    output wire signed [63:0] matmult_out_b69,
    output wire signed [63:0] matmult_out_b70,
    output wire signed [63:0] matmult_out_b71,
    output wire signed [63:0] matmult_out_b72,
    output wire signed [63:0] matmult_out_b73,
    output wire signed [63:0] matmult_out_b74,
    output wire signed [63:0] matmult_out_b75,
    output wire signed [63:0] matmult_out_b76,
    output wire signed [63:0] matmult_out_b77,
    output wire signed [63:0] matmult_out_b78,
    output wire signed [63:0] matmult_out_b79,
    output wire signed [63:0] matmult_out_b80,
    output wire signed [63:0] matmult_out_b81,
    output wire signed [63:0] matmult_out_b82,
    output wire signed [63:0] matmult_out_b83,
    output wire signed [63:0] matmult_out_b84,
    output wire signed [63:0] matmult_out_b85,
    output wire signed [63:0] matmult_out_b86,
    output wire signed [63:0] matmult_out_b87,
    output wire signed [63:0] matmult_out_b88,
    output wire signed [63:0] matmult_out_b89,
    output wire signed [63:0] matmult_out_b90,
    output wire signed [63:0] matmult_out_b91,
    output wire signed [63:0] matmult_out_b92,
    output wire signed [63:0] matmult_out_b93,
    output wire signed [63:0] matmult_out_b94,
    output wire signed [63:0] matmult_out_b95,
    output wire signed [63:0] matmult_out_b96,
    output wire signed [63:0] matmult_out_b97,
    output wire signed [63:0] matmult_out_b98,
    output wire signed [63:0] matmult_out_b99,
    output wire signed [63:0] matmult_out_b100,
    output wire signed [63:0] matmult_out_b101,
    output wire signed [63:0] matmult_out_b102,
    output wire signed [63:0] matmult_out_b103,
    output wire signed [63:0] matmult_out_b104,
    output wire signed [63:0] matmult_out_b105,
    output wire signed [63:0] matmult_out_b106,
    output wire signed [63:0] matmult_out_b107,
    output wire signed [63:0] matmult_out_b108,
    output wire signed [63:0] matmult_out_b109,
    output wire signed [63:0] matmult_out_b110,
    output wire signed [63:0] matmult_out_b111,
    output wire signed [63:0] matmult_out_b112,
    output wire signed [63:0] matmult_out_b113,
    output wire signed [63:0] matmult_out_b114,
    output wire signed [63:0] matmult_out_b115,
    output wire signed [63:0] matmult_out_b116,
    output wire signed [63:0] matmult_out_b117,
    output wire signed [63:0] matmult_out_b118,
    output wire signed [63:0] matmult_out_b119,
    output wire signed [63:0] matmult_out_b120,
    output wire signed [63:0] matmult_out_b121,
    output wire signed [63:0] matmult_out_b122,
    output wire signed [63:0] matmult_out_b123,
    output wire signed [63:0] matmult_out_b124,
    output wire signed [63:0] matmult_out_b125,
    output wire signed [63:0] matmult_out_b126,
    output wire signed [63:0] matmult_out_b127,
    output wire signed [63:0] matmult_out_b128,
    output wire signed [63:0] matmult_out_b129,
    output wire signed [63:0] matmult_out_b130,
    output wire signed [63:0] matmult_out_b131,
    output wire signed [63:0] matmult_out_b132,
    output wire signed [63:0] matmult_out_b133,
    output wire signed [63:0] matmult_out_b134,
    output wire signed [63:0] matmult_out_b135,
    output wire signed [63:0] matmult_out_b136,
    output wire signed [63:0] matmult_out_b137,
    output wire signed [63:0] matmult_out_b138,
    output wire signed [63:0] matmult_out_b139,
    output wire signed [63:0] matmult_out_b140,
    output wire signed [63:0] matmult_out_b141,
    output wire signed [63:0] matmult_out_b142,
    output wire signed [63:0] matmult_out_b143,
    output wire signed [63:0] matmult_out_b144,
    output wire signed [63:0] matmult_out_b145,
    output wire signed [63:0] matmult_out_b146,
    output wire signed [63:0] matmult_out_b147,
    output wire signed [63:0] matmult_out_b148,
    output wire signed [63:0] matmult_out_b149,
    output wire signed [63:0] matmult_out_b150,
    output wire signed [63:0] matmult_out_b151,
    output wire signed [63:0] matmult_out_b152,
    output wire signed [63:0] matmult_out_b153,
    output wire signed [63:0] matmult_out_b154,
    output wire signed [63:0] matmult_out_b155,
    output wire signed [63:0] matmult_out_b156,
    output wire signed [63:0] matmult_out_b157,
    output wire signed [63:0] matmult_out_b158,
    output wire signed [63:0] matmult_out_b159,
    output wire signed [63:0] matmult_out_b160,
    output wire signed [63:0] matmult_out_b161,
    output wire signed [63:0] matmult_out_b162,
    output wire signed [63:0] matmult_out_b163,
    output wire signed [63:0] matmult_out_b164,
    output wire signed [63:0] matmult_out_b165,
    output wire signed [63:0] matmult_out_b166,
    output wire signed [63:0] matmult_out_b167,
    output wire signed [63:0] matmult_out_b168,
    output wire signed [63:0] matmult_out_b169,
    output wire signed [63:0] matmult_out_b170,
    output wire signed [63:0] matmult_out_b171,
    output wire signed [63:0] matmult_out_b172,
    output wire signed [63:0] matmult_out_b173,
    output wire signed [63:0] matmult_out_b174,
    output wire signed [63:0] matmult_out_b175,
    output wire signed [63:0] matmult_out_b176,
    output wire signed [63:0] matmult_out_b177,
    output wire signed [63:0] matmult_out_b178,
    output wire signed [63:0] matmult_out_b179,
    output wire signed [63:0] matmult_out_b180,
    output wire signed [63:0] matmult_out_b181,
    output wire signed [63:0] matmult_out_b182,
    output wire signed [63:0] matmult_out_b183,
    output wire signed [63:0] matmult_out_b184,
    output wire signed [63:0] matmult_out_b185,
    output wire signed [63:0] matmult_out_b186,
    output wire signed [63:0] matmult_out_b187,
    output wire signed [63:0] matmult_out_b188,
    output wire signed [63:0] matmult_out_b189,
    output wire signed [63:0] matmult_out_b190,
    output wire signed [63:0] matmult_out_b191,
    output wire signed [63:0] matmult_out_b192,
    output wire signed [63:0] matmult_out_b193,
    output wire signed [63:0] matmult_out_b194,
    output wire signed [63:0] matmult_out_b195,
    output wire signed [63:0] matmult_out_b196,
    output wire signed [63:0] matmult_out_b197,
    output wire signed [63:0] matmult_out_b198,
    output wire signed [63:0] matmult_out_b199,
    output wire signed [63:0] matmult_out_b200,
    output wire signed [63:0] matmult_out_b201,
    output wire signed [63:0] matmult_out_b202,
    output wire signed [63:0] matmult_out_b203,
    output wire signed [63:0] matmult_out_b204,
    output wire signed [63:0] matmult_out_b205,
    output wire signed [63:0] matmult_out_b206,
    output wire signed [63:0] matmult_out_b207,
    output wire signed [63:0] matmult_out_b208,
    output wire signed [63:0] matmult_out_b209,
    output wire signed [63:0] matmult_out_b210,
    output wire signed [63:0] matmult_out_b211,
    output wire signed [63:0] matmult_out_b212,
    output wire signed [63:0] matmult_out_b213,
    output wire signed [63:0] matmult_out_b214,
    output wire signed [63:0] matmult_out_b215,
    output wire signed [63:0] matmult_out_b216,
    output wire signed [63:0] matmult_out_b217,
    output wire signed [63:0] matmult_out_b218,
    output wire signed [63:0] matmult_out_b219,
    output wire signed [63:0] matmult_out_b220,
    output wire signed [63:0] matmult_out_b221,
    output wire signed [63:0] matmult_out_b222,
    output wire signed [63:0] matmult_out_b223,
    output wire signed [63:0] matmult_out_b224,
    output wire signed [63:0] matmult_out_b225,
    output wire signed [63:0] matmult_out_b226,
    output wire signed [63:0] matmult_out_b227,
    output wire signed [63:0] matmult_out_b228,
    output wire signed [63:0] matmult_out_b229,
    output wire signed [63:0] matmult_out_b230,
    output wire signed [63:0] matmult_out_b231,
    output wire signed [63:0] matmult_out_b232,
    output wire signed [63:0] matmult_out_b233,
    output wire signed [63:0] matmult_out_b234,
    output wire signed [63:0] matmult_out_b235,
    output wire signed [63:0] matmult_out_b236,
    output wire signed [63:0] matmult_out_b237,
    output wire signed [63:0] matmult_out_b238,
    output wire signed [63:0] matmult_out_b239,
    output wire signed [63:0] matmult_out_b240,
    output wire signed [63:0] matmult_out_b241,
    output wire signed [63:0] matmult_out_b242,
    output wire signed [63:0] matmult_out_b243,
    output wire signed [63:0] matmult_out_b244,
    output wire signed [63:0] matmult_out_b245,
    output wire signed [63:0] matmult_out_b246,
    output wire signed [63:0] matmult_out_b247,
    output wire signed [63:0] matmult_out_b248,
    output wire signed [63:0] matmult_out_b249,
    output wire signed [63:0] matmult_out_b250,
    output wire signed [63:0] matmult_out_b251,
    output wire signed [63:0] matmult_out_b252,
    output wire signed [63:0] matmult_out_b253,
    output wire signed [63:0] matmult_out_b254,
    output wire signed [63:0] matmult_out_b255,
    output wire signed [63:0] matmult_out_b256,
    output wire signed [63:0] matmult_out_b257,
    output wire signed [63:0] matmult_out_b258,
    output wire signed [63:0] matmult_out_b259,
    output wire signed [63:0] matmult_out_b260,
    output wire signed [63:0] matmult_out_b261,
    output wire signed [63:0] matmult_out_b262,
    output wire signed [63:0] matmult_out_b263,
    output wire signed [63:0] matmult_out_b264,
    output wire signed [63:0] matmult_out_b265,
    output wire signed [63:0] matmult_out_b266,
    output wire signed [63:0] matmult_out_b267,
    output wire signed [63:0] matmult_out_b268,
    output wire signed [63:0] matmult_out_b269,
    output wire signed [63:0] matmult_out_b270,
    output wire signed [63:0] matmult_out_b271,
    output wire signed [63:0] matmult_out_b272,
    output wire signed [63:0] matmult_out_b273,
    output wire signed [63:0] matmult_out_b274,
    output wire signed [63:0] matmult_out_b275,
    output wire signed [63:0] matmult_out_b276,
    output wire signed [63:0] matmult_out_b277,
    output wire signed [63:0] matmult_out_b278,
    output wire signed [63:0] matmult_out_b279,
    input wire [7:0] matmult_in_col,
    input wire signed [63:0] matmult_in_c0,
    input wire signed [63:0] matmult_in_c1,
    input wire signed [63:0] matmult_in_c2,
    input wire signed [63:0] matmult_in_c3,
    input wire signed [63:0] matmult_in_c4,
    input wire signed [63:0] matmult_in_c5,
    input wire signed [63:0] matmult_in_c6,
    input wire signed [63:0] matmult_in_c7,
    input wire signed [63:0] matmult_in_c8,
    input wire signed [63:0] matmult_in_c9,
    input wire signed [63:0] matmult_in_c10,
    input wire signed [63:0] matmult_in_c11,
    input wire signed [63:0] matmult_in_c12,
    input wire signed [63:0] matmult_in_c13,
    input wire signed [63:0] matmult_in_c14,
    input wire signed [63:0] matmult_in_c15,
    input wire signed [63:0] matmult_in_c16,
    input wire signed [63:0] matmult_in_c17,
    input wire signed [63:0] matmult_in_c18,
    input wire signed [63:0] matmult_in_c19,
    input wire signed [63:0] matmult_in_c20,
    input wire signed [63:0] matmult_in_c21,
    input wire signed [63:0] matmult_in_c22,
    input wire signed [63:0] matmult_in_c23,
    input wire signed [63:0] matmult_in_c24,
    input wire signed [63:0] matmult_in_c25,
    input wire signed [63:0] matmult_in_c26,
    input wire signed [63:0] matmult_in_c27,
    input wire signed [63:0] matmult_in_c28,
    input wire signed [63:0] matmult_in_c29,
    input wire signed [63:0] matmult_in_c30,
    input wire signed [63:0] matmult_in_c31,
    input wire signed [63:0] matmult_in_c32,
    input wire signed [63:0] matmult_in_c33,
    input wire signed [63:0] matmult_in_c34,
    input wire signed [63:0] matmult_in_c35,
    input wire signed [63:0] matmult_in_c36,
    input wire signed [63:0] matmult_in_c37,
    input wire signed [63:0] matmult_in_c38,
    input wire signed [63:0] matmult_in_c39,
    input wire signed [63:0] matmult_in_c40,
    input wire signed [63:0] matmult_in_c41,
    input wire signed [63:0] matmult_in_c42,
    input wire signed [63:0] matmult_in_c43,
    input wire signed [63:0] matmult_in_c44,
    input wire signed [63:0] matmult_in_c45,
    input wire signed [63:0] matmult_in_c46,
    input wire signed [63:0] matmult_in_c47,
    input wire signed [63:0] matmult_in_c48,
    input wire signed [63:0] matmult_in_c49,
    input wire signed [63:0] matmult_in_c50,
    input wire signed [63:0] matmult_in_c51,
    input wire signed [63:0] matmult_in_c52,
    input wire signed [63:0] matmult_in_c53,
    input wire signed [63:0] matmult_in_c54,
    input wire signed [63:0] matmult_in_c55,
    input wire signed [63:0] matmult_in_c56,
    input wire signed [63:0] matmult_in_c57,
    input wire signed [63:0] matmult_in_c58,
    input wire signed [63:0] matmult_in_c59,
    input wire signed [63:0] matmult_in_c60,
    input wire signed [63:0] matmult_in_c61,
    input wire signed [63:0] matmult_in_c62,
    input wire signed [63:0] matmult_in_c63,
    input wire signed [63:0] matmult_in_c64,
    input wire signed [63:0] matmult_in_c65,
    input wire signed [63:0] matmult_in_c66,
    input wire signed [63:0] matmult_in_c67,
    input wire signed [63:0] matmult_in_c68,
    input wire signed [63:0] matmult_in_c69,
    input wire signed [63:0] matmult_in_c70,
    input wire signed [63:0] matmult_in_c71,
    input wire signed [63:0] matmult_in_c72,
    input wire signed [63:0] matmult_in_c73,
    input wire signed [63:0] matmult_in_c74,
    input wire signed [63:0] matmult_in_c75,
    input wire signed [63:0] matmult_in_c76,
    input wire signed [63:0] matmult_in_c77,
    input wire signed [63:0] matmult_in_c78,
    input wire signed [63:0] matmult_in_c79,
    input wire signed [63:0] matmult_in_c80,
    input wire signed [63:0] matmult_in_c81,
    input wire signed [63:0] matmult_in_c82,
    input wire signed [63:0] matmult_in_c83,
    input wire signed [63:0] matmult_in_c84,
    input wire signed [63:0] matmult_in_c85,
    input wire signed [63:0] matmult_in_c86,
    input wire signed [63:0] matmult_in_c87,
    input wire signed [63:0] matmult_in_c88,
    input wire signed [63:0] matmult_in_c89,
    input wire signed [63:0] matmult_in_c90,
    input wire signed [63:0] matmult_in_c91,
    input wire signed [63:0] matmult_in_c92,
    input wire signed [63:0] matmult_in_c93,
    input wire signed [63:0] matmult_in_c94,
    input wire signed [63:0] matmult_in_c95,
    input wire signed [63:0] matmult_in_c96,
    input wire signed [63:0] matmult_in_c97,
    input wire signed [63:0] matmult_in_c98,
    input wire signed [63:0] matmult_in_c99,
    input wire signed [63:0] matmult_in_c100,
    input wire signed [63:0] matmult_in_c101,
    input wire signed [63:0] matmult_in_c102,
    input wire signed [63:0] matmult_in_c103,
    input wire signed [63:0] matmult_in_c104,
    input wire signed [63:0] matmult_in_c105,
    input wire signed [63:0] matmult_in_c106,
    input wire signed [63:0] matmult_in_c107,
    input wire signed [63:0] matmult_in_c108,
    input wire signed [63:0] matmult_in_c109,
    input wire signed [63:0] matmult_in_c110,
    input wire signed [63:0] matmult_in_c111,
    input wire signed [63:0] matmult_in_c112,
    input wire signed [63:0] matmult_in_c113,
    input wire signed [63:0] matmult_in_c114,
    input wire signed [63:0] matmult_in_c115,
    input wire signed [63:0] matmult_in_c116,
    input wire signed [63:0] matmult_in_c117,
    input wire signed [63:0] matmult_in_c118,
    input wire signed [63:0] matmult_in_c119,
    input wire signed [63:0] matmult_in_c120,
    input wire signed [63:0] matmult_in_c121,
    input wire signed [63:0] matmult_in_c122,
    input wire signed [63:0] matmult_in_c123,
    input wire signed [63:0] matmult_in_c124,
    input wire signed [63:0] matmult_in_c125,
    input wire signed [63:0] matmult_in_c126,
    input wire signed [63:0] matmult_in_c127,
    input wire signed [63:0] matmult_in_c128,
    input wire signed [63:0] matmult_in_c129,
    input wire signed [63:0] matmult_in_c130,
    input wire signed [63:0] matmult_in_c131,
    input wire signed [63:0] matmult_in_c132,
    input wire signed [63:0] matmult_in_c133,
    input wire signed [63:0] matmult_in_c134,
    input wire signed [63:0] matmult_in_c135,
    input wire signed [63:0] matmult_in_c136,
    input wire signed [63:0] matmult_in_c137,
    input wire signed [63:0] matmult_in_c138,
    input wire signed [63:0] matmult_in_c139,
    input wire signed [63:0] matmult_in_c140,
    input wire signed [63:0] matmult_in_c141,
    input wire signed [63:0] matmult_in_c142,
    input wire signed [63:0] matmult_in_c143,
    input wire signed [63:0] matmult_in_c144,
    input wire signed [63:0] matmult_in_c145,
    input wire signed [63:0] matmult_in_c146,
    input wire signed [63:0] matmult_in_c147,
    input wire signed [63:0] matmult_in_c148,
    input wire signed [63:0] matmult_in_c149,
    input wire signed [63:0] matmult_in_c150,
    input wire signed [63:0] matmult_in_c151,
    input wire signed [63:0] matmult_in_c152,
    input wire signed [63:0] matmult_in_c153,
    input wire signed [63:0] matmult_in_c154,
    input wire signed [63:0] matmult_in_c155,
    input wire signed [63:0] matmult_in_c156,
    input wire signed [63:0] matmult_in_c157,
    input wire signed [63:0] matmult_in_c158,
    input wire signed [63:0] matmult_in_c159,
    input wire signed [63:0] matmult_in_c160,
    input wire signed [63:0] matmult_in_c161,
    input wire signed [63:0] matmult_in_c162,
    input wire signed [63:0] matmult_in_c163,
    input wire signed [63:0] matmult_in_c164,
    input wire signed [63:0] matmult_in_c165,
    input wire signed [63:0] matmult_in_c166,
    input wire signed [63:0] matmult_in_c167,
    input wire signed [63:0] matmult_in_c168,
    input wire signed [63:0] matmult_in_c169,
    input wire signed [63:0] matmult_in_c170,
    input wire signed [63:0] matmult_in_c171,
    input wire signed [63:0] matmult_in_c172,
    input wire signed [63:0] matmult_in_c173,
    input wire signed [63:0] matmult_in_c174,
    input wire signed [63:0] matmult_in_c175,
    input wire signed [63:0] matmult_in_c176,
    input wire signed [63:0] matmult_in_c177,
    input wire signed [63:0] matmult_in_c178,
    input wire signed [63:0] matmult_in_c179,
    input wire signed [63:0] matmult_in_c180,
    input wire signed [63:0] matmult_in_c181,
    input wire signed [63:0] matmult_in_c182,
    input wire signed [63:0] matmult_in_c183,
    input wire signed [63:0] matmult_in_c184,
    input wire signed [63:0] matmult_in_c185,
    input wire signed [63:0] matmult_in_c186,
    input wire signed [63:0] matmult_in_c187,
    input wire signed [63:0] matmult_in_c188,
    input wire signed [63:0] matmult_in_c189,
    input wire signed [63:0] matmult_in_c190,
    input wire signed [63:0] matmult_in_c191,
    input wire signed [63:0] matmult_in_c192,
    input wire signed [63:0] matmult_in_c193,
    input wire signed [63:0] matmult_in_c194,
    input wire signed [63:0] matmult_in_c195,
    input wire signed [63:0] matmult_in_c196,
    input wire signed [63:0] matmult_in_c197,
    input wire signed [63:0] matmult_in_c198,
    input wire signed [63:0] matmult_in_c199,
    input wire signed [63:0] matmult_in_c200,
    input wire signed [63:0] matmult_in_c201,
    input wire signed [63:0] matmult_in_c202,
    input wire signed [63:0] matmult_in_c203,
    input wire signed [63:0] matmult_in_c204,
    input wire signed [63:0] matmult_in_c205,
    input wire signed [63:0] matmult_in_c206,
    input wire signed [63:0] matmult_in_c207,
    input wire signed [63:0] matmult_in_c208,
    input wire signed [63:0] matmult_in_c209,
    input wire signed [63:0] matmult_in_c210,
    input wire signed [63:0] matmult_in_c211,
    input wire signed [63:0] matmult_in_c212,
    input wire signed [63:0] matmult_in_c213,
    input wire signed [63:0] matmult_in_c214,
    input wire signed [63:0] matmult_in_c215,
    input wire signed [63:0] matmult_in_c216,
    input wire signed [63:0] matmult_in_c217,
    input wire signed [63:0] matmult_in_c218,
    input wire signed [63:0] matmult_in_c219,
    input wire signed [63:0] matmult_in_c220,
    input wire signed [63:0] matmult_in_c221,
    input wire signed [63:0] matmult_in_c222,
    input wire signed [63:0] matmult_in_c223,
    input wire signed [63:0] matmult_in_c224,
    input wire signed [63:0] matmult_in_c225,
    input wire signed [63:0] matmult_in_c226,
    input wire signed [63:0] matmult_in_c227,
    input wire signed [63:0] matmult_in_c228,
    input wire signed [63:0] matmult_in_c229,
    input wire signed [63:0] matmult_in_c230,
    input wire signed [63:0] matmult_in_c231,
    input wire signed [63:0] matmult_in_c232,
    input wire signed [63:0] matmult_in_c233,
    input wire signed [63:0] matmult_in_c234,
    input wire signed [63:0] matmult_in_c235,
    input wire signed [63:0] matmult_in_c236,
    input wire signed [63:0] matmult_in_c237,
    input wire signed [63:0] matmult_in_c238,
    input wire signed [63:0] matmult_in_c239,
    input wire signed [63:0] matmult_in_c240,
    input wire signed [63:0] matmult_in_c241,
    input wire signed [63:0] matmult_in_c242,
    input wire signed [63:0] matmult_in_c243,
    input wire signed [63:0] matmult_in_c244,
    input wire signed [63:0] matmult_in_c245,
    input wire signed [63:0] matmult_in_c246,
    input wire signed [63:0] matmult_in_c247,
    input wire signed [63:0] matmult_in_c248,
    input wire signed [63:0] matmult_in_c249,
    input wire signed [63:0] matmult_in_c250,
    input wire signed [63:0] matmult_in_c251,
    input wire signed [63:0] matmult_in_c252,
    input wire signed [63:0] matmult_in_c253,
    input wire signed [63:0] matmult_in_c254,
    input wire signed [63:0] matmult_in_c255,
    input wire signed [63:0] matmult_in_c256,
    input wire signed [63:0] matmult_in_c257,
    input wire signed [63:0] matmult_in_c258,
    input wire signed [63:0] matmult_in_c259,
    input wire signed [63:0] matmult_in_c260,
    input wire signed [63:0] matmult_in_c261,
    input wire signed [63:0] matmult_in_c262,
    input wire signed [63:0] matmult_in_c263,
    input wire signed [63:0] matmult_in_c264,
    input wire signed [63:0] matmult_in_c265,
    input wire signed [63:0] matmult_in_c266,
    input wire signed [63:0] matmult_in_c267,
    input wire signed [63:0] matmult_in_c268,
    input wire signed [63:0] matmult_in_c269,
    input wire signed [63:0] matmult_in_c270,
    input wire signed [63:0] matmult_in_c271,
    input wire signed [63:0] matmult_in_c272,
    input wire signed [63:0] matmult_in_c273,
    input wire signed [63:0] matmult_in_c274,
    input wire signed [63:0] matmult_in_c275,
    input wire signed [63:0] matmult_in_c276,
    input wire signed [63:0] matmult_in_c277,
    input wire signed [63:0] matmult_in_c278,
    input wire signed [63:0] matmult_in_c279,
    output wire signed [63:0] matmult_out_c0,
    output wire signed [63:0] matmult_out_c1,
    output wire signed [63:0] matmult_out_c2,
    output wire signed [63:0] matmult_out_c3,
    output wire signed [63:0] matmult_out_c4,
    output wire signed [63:0] matmult_out_c5,
    output wire signed [63:0] matmult_out_c6,
    output wire signed [63:0] matmult_out_c7,
    output wire signed [63:0] matmult_out_c8,
    output wire signed [63:0] matmult_out_c9,
    output wire signed [63:0] matmult_out_c10,
    output wire signed [63:0] matmult_out_c11,
    output wire signed [63:0] matmult_out_c12,
    output wire signed [63:0] matmult_out_c13,
    output wire signed [63:0] matmult_out_c14,
    output wire signed [63:0] matmult_out_c15,
    output wire signed [63:0] matmult_out_c16,
    output wire signed [63:0] matmult_out_c17,
    output wire signed [63:0] matmult_out_c18,
    output wire signed [63:0] matmult_out_c19,
    output wire signed [63:0] matmult_out_c20,
    output wire signed [63:0] matmult_out_c21,
    output wire signed [63:0] matmult_out_c22,
    output wire signed [63:0] matmult_out_c23,
    output wire signed [63:0] matmult_out_c24,
    output wire signed [63:0] matmult_out_c25,
    output wire signed [63:0] matmult_out_c26,
    output wire signed [63:0] matmult_out_c27,
    output wire signed [63:0] matmult_out_c28,
    output wire signed [63:0] matmult_out_c29,
    output wire signed [63:0] matmult_out_c30,
    output wire signed [63:0] matmult_out_c31,
    output wire signed [63:0] matmult_out_c32,
    output wire signed [63:0] matmult_out_c33,
    output wire signed [63:0] matmult_out_c34,
    output wire signed [63:0] matmult_out_c35,
    output wire signed [63:0] matmult_out_c36,
    output wire signed [63:0] matmult_out_c37,
    output wire signed [63:0] matmult_out_c38,
    output wire signed [63:0] matmult_out_c39,
    output wire signed [63:0] matmult_out_c40,
    output wire signed [63:0] matmult_out_c41,
    output wire signed [63:0] matmult_out_c42,
    output wire signed [63:0] matmult_out_c43,
    output wire signed [63:0] matmult_out_c44,
    output wire signed [63:0] matmult_out_c45,
    output wire signed [63:0] matmult_out_c46,
    output wire signed [63:0] matmult_out_c47,
    output wire signed [63:0] matmult_out_c48,
    output wire signed [63:0] matmult_out_c49,
    output wire signed [63:0] matmult_out_c50,
    output wire signed [63:0] matmult_out_c51,
    output wire signed [63:0] matmult_out_c52,
    output wire signed [63:0] matmult_out_c53,
    output wire signed [63:0] matmult_out_c54,
    output wire signed [63:0] matmult_out_c55,
    output wire signed [63:0] matmult_out_c56,
    output wire signed [63:0] matmult_out_c57,
    output wire signed [63:0] matmult_out_c58,
    output wire signed [63:0] matmult_out_c59,
    output wire signed [63:0] matmult_out_c60,
    output wire signed [63:0] matmult_out_c61,
    output wire signed [63:0] matmult_out_c62,
    output wire signed [63:0] matmult_out_c63,
    output wire signed [63:0] matmult_out_c64,
    output wire signed [63:0] matmult_out_c65,
    output wire signed [63:0] matmult_out_c66,
    output wire signed [63:0] matmult_out_c67,
    output wire signed [63:0] matmult_out_c68,
    output wire signed [63:0] matmult_out_c69,
    output wire signed [63:0] matmult_out_c70,
    output wire signed [63:0] matmult_out_c71,
    output wire signed [63:0] matmult_out_c72,
    output wire signed [63:0] matmult_out_c73,
    output wire signed [63:0] matmult_out_c74,
    output wire signed [63:0] matmult_out_c75,
    output wire signed [63:0] matmult_out_c76,
    output wire signed [63:0] matmult_out_c77,
    output wire signed [63:0] matmult_out_c78,
    output wire signed [63:0] matmult_out_c79,
    output wire signed [63:0] matmult_out_c80,
    output wire signed [63:0] matmult_out_c81,
    output wire signed [63:0] matmult_out_c82,
    output wire signed [63:0] matmult_out_c83,
    output wire signed [63:0] matmult_out_c84,
    output wire signed [63:0] matmult_out_c85,
    output wire signed [63:0] matmult_out_c86,
    output wire signed [63:0] matmult_out_c87,
    output wire signed [63:0] matmult_out_c88,
    output wire signed [63:0] matmult_out_c89,
    output wire signed [63:0] matmult_out_c90,
    output wire signed [63:0] matmult_out_c91,
    output wire signed [63:0] matmult_out_c92,
    output wire signed [63:0] matmult_out_c93,
    output wire signed [63:0] matmult_out_c94,
    output wire signed [63:0] matmult_out_c95,
    output wire signed [63:0] matmult_out_c96,
    output wire signed [63:0] matmult_out_c97,
    output wire signed [63:0] matmult_out_c98,
    output wire signed [63:0] matmult_out_c99,
    output wire signed [63:0] matmult_out_c100,
    output wire signed [63:0] matmult_out_c101,
    output wire signed [63:0] matmult_out_c102,
    output wire signed [63:0] matmult_out_c103,
    output wire signed [63:0] matmult_out_c104,
    output wire signed [63:0] matmult_out_c105,
    output wire signed [63:0] matmult_out_c106,
    output wire signed [63:0] matmult_out_c107,
    output wire signed [63:0] matmult_out_c108,
    output wire signed [63:0] matmult_out_c109,
    output wire signed [63:0] matmult_out_c110,
    output wire signed [63:0] matmult_out_c111,
    output wire signed [63:0] matmult_out_c112,
    output wire signed [63:0] matmult_out_c113,
    output wire signed [63:0] matmult_out_c114,
    output wire signed [63:0] matmult_out_c115,
    output wire signed [63:0] matmult_out_c116,
    output wire signed [63:0] matmult_out_c117,
    output wire signed [63:0] matmult_out_c118,
    output wire signed [63:0] matmult_out_c119,
    output wire signed [63:0] matmult_out_c120,
    output wire signed [63:0] matmult_out_c121,
    output wire signed [63:0] matmult_out_c122,
    output wire signed [63:0] matmult_out_c123,
    output wire signed [63:0] matmult_out_c124,
    output wire signed [63:0] matmult_out_c125,
    output wire signed [63:0] matmult_out_c126,
    output wire signed [63:0] matmult_out_c127,
    output wire signed [63:0] matmult_out_c128,
    output wire signed [63:0] matmult_out_c129,
    output wire signed [63:0] matmult_out_c130,
    output wire signed [63:0] matmult_out_c131,
    output wire signed [63:0] matmult_out_c132,
    output wire signed [63:0] matmult_out_c133,
    output wire signed [63:0] matmult_out_c134,
    output wire signed [63:0] matmult_out_c135,
    output wire signed [63:0] matmult_out_c136,
    output wire signed [63:0] matmult_out_c137,
    output wire signed [63:0] matmult_out_c138,
    output wire signed [63:0] matmult_out_c139,
    output wire signed [63:0] matmult_out_c140,
    output wire signed [63:0] matmult_out_c141,
    output wire signed [63:0] matmult_out_c142,
    output wire signed [63:0] matmult_out_c143,
    output wire signed [63:0] matmult_out_c144,
    output wire signed [63:0] matmult_out_c145,
    output wire signed [63:0] matmult_out_c146,
    output wire signed [63:0] matmult_out_c147,
    output wire signed [63:0] matmult_out_c148,
    output wire signed [63:0] matmult_out_c149,
    output wire signed [63:0] matmult_out_c150,
    output wire signed [63:0] matmult_out_c151,
    output wire signed [63:0] matmult_out_c152,
    output wire signed [63:0] matmult_out_c153,
    output wire signed [63:0] matmult_out_c154,
    output wire signed [63:0] matmult_out_c155,
    output wire signed [63:0] matmult_out_c156,
    output wire signed [63:0] matmult_out_c157,
    output wire signed [63:0] matmult_out_c158,
    output wire signed [63:0] matmult_out_c159,
    output wire signed [63:0] matmult_out_c160,
    output wire signed [63:0] matmult_out_c161,
    output wire signed [63:0] matmult_out_c162,
    output wire signed [63:0] matmult_out_c163,
    output wire signed [63:0] matmult_out_c164,
    output wire signed [63:0] matmult_out_c165,
    output wire signed [63:0] matmult_out_c166,
    output wire signed [63:0] matmult_out_c167,
    output wire signed [63:0] matmult_out_c168,
    output wire signed [63:0] matmult_out_c169,
    output wire signed [63:0] matmult_out_c170,
    output wire signed [63:0] matmult_out_c171,
    output wire signed [63:0] matmult_out_c172,
    output wire signed [63:0] matmult_out_c173,
    output wire signed [63:0] matmult_out_c174,
    output wire signed [63:0] matmult_out_c175,
    output wire signed [63:0] matmult_out_c176,
    output wire signed [63:0] matmult_out_c177,
    output wire signed [63:0] matmult_out_c178,
    output wire signed [63:0] matmult_out_c179,
    output wire signed [63:0] matmult_out_c180,
    output wire signed [63:0] matmult_out_c181,
    output wire signed [63:0] matmult_out_c182,
    output wire signed [63:0] matmult_out_c183,
    output wire signed [63:0] matmult_out_c184,
    output wire signed [63:0] matmult_out_c185,
    output wire signed [63:0] matmult_out_c186,
    output wire signed [63:0] matmult_out_c187,
    output wire signed [63:0] matmult_out_c188,
    output wire signed [63:0] matmult_out_c189,
    output wire signed [63:0] matmult_out_c190,
    output wire signed [63:0] matmult_out_c191,
    output wire signed [63:0] matmult_out_c192,
    output wire signed [63:0] matmult_out_c193,
    output wire signed [63:0] matmult_out_c194,
    output wire signed [63:0] matmult_out_c195,
    output wire signed [63:0] matmult_out_c196,
    output wire signed [63:0] matmult_out_c197,
    output wire signed [63:0] matmult_out_c198,
    output wire signed [63:0] matmult_out_c199,
    output wire signed [63:0] matmult_out_c200,
    output wire signed [63:0] matmult_out_c201,
    output wire signed [63:0] matmult_out_c202,
    output wire signed [63:0] matmult_out_c203,
    output wire signed [63:0] matmult_out_c204,
    output wire signed [63:0] matmult_out_c205,
    output wire signed [63:0] matmult_out_c206,
    output wire signed [63:0] matmult_out_c207,
    output wire signed [63:0] matmult_out_c208,
    output wire signed [63:0] matmult_out_c209,
    output wire signed [63:0] matmult_out_c210,
    output wire signed [63:0] matmult_out_c211,
    output wire signed [63:0] matmult_out_c212,
    output wire signed [63:0] matmult_out_c213,
    output wire signed [63:0] matmult_out_c214,
    output wire signed [63:0] matmult_out_c215,
    output wire signed [63:0] matmult_out_c216,
    output wire signed [63:0] matmult_out_c217,
    output wire signed [63:0] matmult_out_c218,
    output wire signed [63:0] matmult_out_c219,
    output wire signed [63:0] matmult_out_c220,
    output wire signed [63:0] matmult_out_c221,
    output wire signed [63:0] matmult_out_c222,
    output wire signed [63:0] matmult_out_c223,
    output wire signed [63:0] matmult_out_c224,
    output wire signed [63:0] matmult_out_c225,
    output wire signed [63:0] matmult_out_c226,
    output wire signed [63:0] matmult_out_c227,
    output wire signed [63:0] matmult_out_c228,
    output wire signed [63:0] matmult_out_c229,
    output wire signed [63:0] matmult_out_c230,
    output wire signed [63:0] matmult_out_c231,
    output wire signed [63:0] matmult_out_c232,
    output wire signed [63:0] matmult_out_c233,
    output wire signed [63:0] matmult_out_c234,
    output wire signed [63:0] matmult_out_c235,
    output wire signed [63:0] matmult_out_c236,
    output wire signed [63:0] matmult_out_c237,
    output wire signed [63:0] matmult_out_c238,
    output wire signed [63:0] matmult_out_c239,
    output wire signed [63:0] matmult_out_c240,
    output wire signed [63:0] matmult_out_c241,
    output wire signed [63:0] matmult_out_c242,
    output wire signed [63:0] matmult_out_c243,
    output wire signed [63:0] matmult_out_c244,
    output wire signed [63:0] matmult_out_c245,
    output wire signed [63:0] matmult_out_c246,
    output wire signed [63:0] matmult_out_c247,
    output wire signed [63:0] matmult_out_c248,
    output wire signed [63:0] matmult_out_c249,
    output wire signed [63:0] matmult_out_c250,
    output wire signed [63:0] matmult_out_c251,
    output wire signed [63:0] matmult_out_c252,
    output wire signed [63:0] matmult_out_c253,
    output wire signed [63:0] matmult_out_c254,
    output wire signed [63:0] matmult_out_c255,
    output wire signed [63:0] matmult_out_c256,
    output wire signed [63:0] matmult_out_c257,
    output wire signed [63:0] matmult_out_c258,
    output wire signed [63:0] matmult_out_c259,
    output wire signed [63:0] matmult_out_c260,
    output wire signed [63:0] matmult_out_c261,
    output wire signed [63:0] matmult_out_c262,
    output wire signed [63:0] matmult_out_c263,
    output wire signed [63:0] matmult_out_c264,
    output wire signed [63:0] matmult_out_c265,
    output wire signed [63:0] matmult_out_c266,
    output wire signed [63:0] matmult_out_c267,
    output wire signed [63:0] matmult_out_c268,
    output wire signed [63:0] matmult_out_c269,
    output wire signed [63:0] matmult_out_c270,
    output wire signed [63:0] matmult_out_c271,
    output wire signed [63:0] matmult_out_c272,
    output wire signed [63:0] matmult_out_c273,
    output wire signed [63:0] matmult_out_c274,
    output wire signed [63:0] matmult_out_c275,
    output wire signed [63:0] matmult_out_c276,
    output wire signed [63:0] matmult_out_c277,
    output wire signed [63:0] matmult_out_c278,
    output wire signed [63:0] matmult_out_c279
);
    localparam idle = 0;
    localparam fin = 1;
    localparam calc = 2;
    reg [63:0] a[0:279];
    reg [63:0] b[0:279];
    reg [63:0] c[0:279];
    reg [1:0] state;

    assign matmult_out_c0 = c[0];
    assign matmult_out_c1 = c[1];
    assign matmult_out_c2 = c[2];
    assign matmult_out_c3 = c[3];
    assign matmult_out_c4 = c[4];
    assign matmult_out_c5 = c[5];
    assign matmult_out_c6 = c[6];
    assign matmult_out_c7 = c[7];
    assign matmult_out_c8 = c[8];
    assign matmult_out_c9 = c[9];
    assign matmult_out_c10 = c[10];
    assign matmult_out_c11 = c[11];
    assign matmult_out_c12 = c[12];
    assign matmult_out_c13 = c[13];
    assign matmult_out_c14 = c[14];
    assign matmult_out_c15 = c[15];
    assign matmult_out_c16 = c[16];
    assign matmult_out_c17 = c[17];
    assign matmult_out_c18 = c[18];
    assign matmult_out_c19 = c[19];
    assign matmult_out_c20 = c[20];
    assign matmult_out_c21 = c[21];
    assign matmult_out_c22 = c[22];
    assign matmult_out_c23 = c[23];
    assign matmult_out_c24 = c[24];
    assign matmult_out_c25 = c[25];
    assign matmult_out_c26 = c[26];
    assign matmult_out_c27 = c[27];
    assign matmult_out_c28 = c[28];
    assign matmult_out_c29 = c[29];
    assign matmult_out_c30 = c[30];
    assign matmult_out_c31 = c[31];
    assign matmult_out_c32 = c[32];
    assign matmult_out_c33 = c[33];
    assign matmult_out_c34 = c[34];
    assign matmult_out_c35 = c[35];
    assign matmult_out_c36 = c[36];
    assign matmult_out_c37 = c[37];
    assign matmult_out_c38 = c[38];
    assign matmult_out_c39 = c[39];
    assign matmult_out_c40 = c[40];
    assign matmult_out_c41 = c[41];
    assign matmult_out_c42 = c[42];
    assign matmult_out_c43 = c[43];
    assign matmult_out_c44 = c[44];
    assign matmult_out_c45 = c[45];
    assign matmult_out_c46 = c[46];
    assign matmult_out_c47 = c[47];
    assign matmult_out_c48 = c[48];
    assign matmult_out_c49 = c[49];
    assign matmult_out_c50 = c[50];
    assign matmult_out_c51 = c[51];
    assign matmult_out_c52 = c[52];
    assign matmult_out_c53 = c[53];
    assign matmult_out_c54 = c[54];
    assign matmult_out_c55 = c[55];
    assign matmult_out_c56 = c[56];
    assign matmult_out_c57 = c[57];
    assign matmult_out_c58 = c[58];
    assign matmult_out_c59 = c[59];
    assign matmult_out_c60 = c[60];
    assign matmult_out_c61 = c[61];
    assign matmult_out_c62 = c[62];
    assign matmult_out_c63 = c[63];
    assign matmult_out_c64 = c[64];
    assign matmult_out_c65 = c[65];
    assign matmult_out_c66 = c[66];
    assign matmult_out_c67 = c[67];
    assign matmult_out_c68 = c[68];
    assign matmult_out_c69 = c[69];
    assign matmult_out_c70 = c[70];
    assign matmult_out_c71 = c[71];
    assign matmult_out_c72 = c[72];
    assign matmult_out_c73 = c[73];
    assign matmult_out_c74 = c[74];
    assign matmult_out_c75 = c[75];
    assign matmult_out_c76 = c[76];
    assign matmult_out_c77 = c[77];
    assign matmult_out_c78 = c[78];
    assign matmult_out_c79 = c[79];
    assign matmult_out_c80 = c[80];
    assign matmult_out_c81 = c[81];
    assign matmult_out_c82 = c[82];
    assign matmult_out_c83 = c[83];
    assign matmult_out_c84 = c[84];
    assign matmult_out_c85 = c[85];
    assign matmult_out_c86 = c[86];
    assign matmult_out_c87 = c[87];
    assign matmult_out_c88 = c[88];
    assign matmult_out_c89 = c[89];
    assign matmult_out_c90 = c[90];
    assign matmult_out_c91 = c[91];
    assign matmult_out_c92 = c[92];
    assign matmult_out_c93 = c[93];
    assign matmult_out_c94 = c[94];
    assign matmult_out_c95 = c[95];
    assign matmult_out_c96 = c[96];
    assign matmult_out_c97 = c[97];
    assign matmult_out_c98 = c[98];
    assign matmult_out_c99 = c[99];
    assign matmult_out_c100 = c[100];
    assign matmult_out_c101 = c[101];
    assign matmult_out_c102 = c[102];
    assign matmult_out_c103 = c[103];
    assign matmult_out_c104 = c[104];
    assign matmult_out_c105 = c[105];
    assign matmult_out_c106 = c[106];
    assign matmult_out_c107 = c[107];
    assign matmult_out_c108 = c[108];
    assign matmult_out_c109 = c[109];
    assign matmult_out_c110 = c[110];
    assign matmult_out_c111 = c[111];
    assign matmult_out_c112 = c[112];
    assign matmult_out_c113 = c[113];
    assign matmult_out_c114 = c[114];
    assign matmult_out_c115 = c[115];
    assign matmult_out_c116 = c[116];
    assign matmult_out_c117 = c[117];
    assign matmult_out_c118 = c[118];
    assign matmult_out_c119 = c[119];
    assign matmult_out_c120 = c[120];
    assign matmult_out_c121 = c[121];
    assign matmult_out_c122 = c[122];
    assign matmult_out_c123 = c[123];
    assign matmult_out_c124 = c[124];
    assign matmult_out_c125 = c[125];
    assign matmult_out_c126 = c[126];
    assign matmult_out_c127 = c[127];
    assign matmult_out_c128 = c[128];
    assign matmult_out_c129 = c[129];
    assign matmult_out_c130 = c[130];
    assign matmult_out_c131 = c[131];
    assign matmult_out_c132 = c[132];
    assign matmult_out_c133 = c[133];
    assign matmult_out_c134 = c[134];
    assign matmult_out_c135 = c[135];
    assign matmult_out_c136 = c[136];
    assign matmult_out_c137 = c[137];
    assign matmult_out_c138 = c[138];
    assign matmult_out_c139 = c[139];
    assign matmult_out_c140 = c[140];
    assign matmult_out_c141 = c[141];
    assign matmult_out_c142 = c[142];
    assign matmult_out_c143 = c[143];
    assign matmult_out_c144 = c[144];
    assign matmult_out_c145 = c[145];
    assign matmult_out_c146 = c[146];
    assign matmult_out_c147 = c[147];
    assign matmult_out_c148 = c[148];
    assign matmult_out_c149 = c[149];
    assign matmult_out_c150 = c[150];
    assign matmult_out_c151 = c[151];
    assign matmult_out_c152 = c[152];
    assign matmult_out_c153 = c[153];
    assign matmult_out_c154 = c[154];
    assign matmult_out_c155 = c[155];
    assign matmult_out_c156 = c[156];
    assign matmult_out_c157 = c[157];
    assign matmult_out_c158 = c[158];
    assign matmult_out_c159 = c[159];
    assign matmult_out_c160 = c[160];
    assign matmult_out_c161 = c[161];
    assign matmult_out_c162 = c[162];
    assign matmult_out_c163 = c[163];
    assign matmult_out_c164 = c[164];
    assign matmult_out_c165 = c[165];
    assign matmult_out_c166 = c[166];
    assign matmult_out_c167 = c[167];
    assign matmult_out_c168 = c[168];
    assign matmult_out_c169 = c[169];
    assign matmult_out_c170 = c[170];
    assign matmult_out_c171 = c[171];
    assign matmult_out_c172 = c[172];
    assign matmult_out_c173 = c[173];
    assign matmult_out_c174 = c[174];
    assign matmult_out_c175 = c[175];
    assign matmult_out_c176 = c[176];
    assign matmult_out_c177 = c[177];
    assign matmult_out_c178 = c[178];
    assign matmult_out_c179 = c[179];
    assign matmult_out_c180 = c[180];
    assign matmult_out_c181 = c[181];
    assign matmult_out_c182 = c[182];
    assign matmult_out_c183 = c[183];
    assign matmult_out_c184 = c[184];
    assign matmult_out_c185 = c[185];
    assign matmult_out_c186 = c[186];
    assign matmult_out_c187 = c[187];
    assign matmult_out_c188 = c[188];
    assign matmult_out_c189 = c[189];
    assign matmult_out_c190 = c[190];
    assign matmult_out_c191 = c[191];
    assign matmult_out_c192 = c[192];
    assign matmult_out_c193 = c[193];
    assign matmult_out_c194 = c[194];
    assign matmult_out_c195 = c[195];
    assign matmult_out_c196 = c[196];
    assign matmult_out_c197 = c[197];
    assign matmult_out_c198 = c[198];
    assign matmult_out_c199 = c[199];
    assign matmult_out_c200 = c[200];
    assign matmult_out_c201 = c[201];
    assign matmult_out_c202 = c[202];
    assign matmult_out_c203 = c[203];
    assign matmult_out_c204 = c[204];
    assign matmult_out_c205 = c[205];
    assign matmult_out_c206 = c[206];
    assign matmult_out_c207 = c[207];
    assign matmult_out_c208 = c[208];
    assign matmult_out_c209 = c[209];
    assign matmult_out_c210 = c[210];
    assign matmult_out_c211 = c[211];
    assign matmult_out_c212 = c[212];
    assign matmult_out_c213 = c[213];
    assign matmult_out_c214 = c[214];
    assign matmult_out_c215 = c[215];
    assign matmult_out_c216 = c[216];
    assign matmult_out_c217 = c[217];
    assign matmult_out_c218 = c[218];
    assign matmult_out_c219 = c[219];
    assign matmult_out_c220 = c[220];
    assign matmult_out_c221 = c[221];
    assign matmult_out_c222 = c[222];
    assign matmult_out_c223 = c[223];
    assign matmult_out_c224 = c[224];
    assign matmult_out_c225 = c[225];
    assign matmult_out_c226 = c[226];
    assign matmult_out_c227 = c[227];
    assign matmult_out_c228 = c[228];
    assign matmult_out_c229 = c[229];
    assign matmult_out_c230 = c[230];
    assign matmult_out_c231 = c[231];
    assign matmult_out_c232 = c[232];
    assign matmult_out_c233 = c[233];
    assign matmult_out_c234 = c[234];
    assign matmult_out_c235 = c[235];
    assign matmult_out_c236 = c[236];
    assign matmult_out_c237 = c[237];
    assign matmult_out_c238 = c[238];
    assign matmult_out_c239 = c[239];
    assign matmult_out_c240 = c[240];
    assign matmult_out_c241 = c[241];
    assign matmult_out_c242 = c[242];
    assign matmult_out_c243 = c[243];
    assign matmult_out_c244 = c[244];
    assign matmult_out_c245 = c[245];
    assign matmult_out_c246 = c[246];
    assign matmult_out_c247 = c[247];
    assign matmult_out_c248 = c[248];
    assign matmult_out_c249 = c[249];
    assign matmult_out_c250 = c[250];
    assign matmult_out_c251 = c[251];
    assign matmult_out_c252 = c[252];
    assign matmult_out_c253 = c[253];
    assign matmult_out_c254 = c[254];
    assign matmult_out_c255 = c[255];
    assign matmult_out_c256 = c[256];
    assign matmult_out_c257 = c[257];
    assign matmult_out_c258 = c[258];
    assign matmult_out_c259 = c[259];
    assign matmult_out_c260 = c[260];
    assign matmult_out_c261 = c[261];
    assign matmult_out_c262 = c[262];
    assign matmult_out_c263 = c[263];
    assign matmult_out_c264 = c[264];
    assign matmult_out_c265 = c[265];
    assign matmult_out_c266 = c[266];
    assign matmult_out_c267 = c[267];
    assign matmult_out_c268 = c[268];
    assign matmult_out_c269 = c[269];
    assign matmult_out_c270 = c[270];
    assign matmult_out_c271 = c[271];
    assign matmult_out_c272 = c[272];
    assign matmult_out_c273 = c[273];
    assign matmult_out_c274 = c[274];
    assign matmult_out_c275 = c[275];
    assign matmult_out_c276 = c[276];
    assign matmult_out_c277 = c[277];
    assign matmult_out_c278 = c[278];
    assign matmult_out_c279 = c[279];

    always @(posedge clk) begin
        if (rst) begin
            for (integer i = 0; i < 280; i++) begin
    a[i] <= 0;
end
            for (integer i = 0; i < 280; i++) begin
    b[i] <= 0;
end
            for (integer i = 0; i < 280; i++) begin
    c[i] <= 0;
end
            state <= 0;
            matmult_valid <= 0;
        end else begin
            case (state)
                idle: begin
                    matmult_valid <= 0;
                    if (matmult_ready) begin
    a[0] <= matmult_in_a0;
    a[1] <= matmult_in_a1;
    a[2] <= matmult_in_a2;
    a[3] <= matmult_in_a3;
    a[4] <= matmult_in_a4;
    a[5] <= matmult_in_a5;
    a[6] <= matmult_in_a6;
    a[7] <= matmult_in_a7;
    a[8] <= matmult_in_a8;
    a[9] <= matmult_in_a9;
    a[10] <= matmult_in_a10;
    a[11] <= matmult_in_a11;
    a[12] <= matmult_in_a12;
    a[13] <= matmult_in_a13;
    a[14] <= matmult_in_a14;
    a[15] <= matmult_in_a15;
    a[16] <= matmult_in_a16;
    a[17] <= matmult_in_a17;
    a[18] <= matmult_in_a18;
    a[19] <= matmult_in_a19;
    a[20] <= matmult_in_a20;
    a[21] <= matmult_in_a21;
    a[22] <= matmult_in_a22;
    a[23] <= matmult_in_a23;
    a[24] <= matmult_in_a24;
    a[25] <= matmult_in_a25;
    a[26] <= matmult_in_a26;
    a[27] <= matmult_in_a27;
    a[28] <= matmult_in_a28;
    a[29] <= matmult_in_a29;
    a[30] <= matmult_in_a30;
    a[31] <= matmult_in_a31;
    a[32] <= matmult_in_a32;
    a[33] <= matmult_in_a33;
    a[34] <= matmult_in_a34;
    a[35] <= matmult_in_a35;
    a[36] <= matmult_in_a36;
    a[37] <= matmult_in_a37;
    a[38] <= matmult_in_a38;
    a[39] <= matmult_in_a39;
    a[40] <= matmult_in_a40;
    a[41] <= matmult_in_a41;
    a[42] <= matmult_in_a42;
    a[43] <= matmult_in_a43;
    a[44] <= matmult_in_a44;
    a[45] <= matmult_in_a45;
    a[46] <= matmult_in_a46;
    a[47] <= matmult_in_a47;
    a[48] <= matmult_in_a48;
    a[49] <= matmult_in_a49;
    a[50] <= matmult_in_a50;
    a[51] <= matmult_in_a51;
    a[52] <= matmult_in_a52;
    a[53] <= matmult_in_a53;
    a[54] <= matmult_in_a54;
    a[55] <= matmult_in_a55;
    a[56] <= matmult_in_a56;
    a[57] <= matmult_in_a57;
    a[58] <= matmult_in_a58;
    a[59] <= matmult_in_a59;
    a[60] <= matmult_in_a60;
    a[61] <= matmult_in_a61;
    a[62] <= matmult_in_a62;
    a[63] <= matmult_in_a63;
    a[64] <= matmult_in_a64;
    a[65] <= matmult_in_a65;
    a[66] <= matmult_in_a66;
    a[67] <= matmult_in_a67;
    a[68] <= matmult_in_a68;
    a[69] <= matmult_in_a69;
    a[70] <= matmult_in_a70;
    a[71] <= matmult_in_a71;
    a[72] <= matmult_in_a72;
    a[73] <= matmult_in_a73;
    a[74] <= matmult_in_a74;
    a[75] <= matmult_in_a75;
    a[76] <= matmult_in_a76;
    a[77] <= matmult_in_a77;
    a[78] <= matmult_in_a78;
    a[79] <= matmult_in_a79;
    a[80] <= matmult_in_a80;
    a[81] <= matmult_in_a81;
    a[82] <= matmult_in_a82;
    a[83] <= matmult_in_a83;
    a[84] <= matmult_in_a84;
    a[85] <= matmult_in_a85;
    a[86] <= matmult_in_a86;
    a[87] <= matmult_in_a87;
    a[88] <= matmult_in_a88;
    a[89] <= matmult_in_a89;
    a[90] <= matmult_in_a90;
    a[91] <= matmult_in_a91;
    a[92] <= matmult_in_a92;
    a[93] <= matmult_in_a93;
    a[94] <= matmult_in_a94;
    a[95] <= matmult_in_a95;
    a[96] <= matmult_in_a96;
    a[97] <= matmult_in_a97;
    a[98] <= matmult_in_a98;
    a[99] <= matmult_in_a99;
    a[100] <= matmult_in_a100;
    a[101] <= matmult_in_a101;
    a[102] <= matmult_in_a102;
    a[103] <= matmult_in_a103;
    a[104] <= matmult_in_a104;
    a[105] <= matmult_in_a105;
    a[106] <= matmult_in_a106;
    a[107] <= matmult_in_a107;
    a[108] <= matmult_in_a108;
    a[109] <= matmult_in_a109;
    a[110] <= matmult_in_a110;
    a[111] <= matmult_in_a111;
    a[112] <= matmult_in_a112;
    a[113] <= matmult_in_a113;
    a[114] <= matmult_in_a114;
    a[115] <= matmult_in_a115;
    a[116] <= matmult_in_a116;
    a[117] <= matmult_in_a117;
    a[118] <= matmult_in_a118;
    a[119] <= matmult_in_a119;
    a[120] <= matmult_in_a120;
    a[121] <= matmult_in_a121;
    a[122] <= matmult_in_a122;
    a[123] <= matmult_in_a123;
    a[124] <= matmult_in_a124;
    a[125] <= matmult_in_a125;
    a[126] <= matmult_in_a126;
    a[127] <= matmult_in_a127;
    a[128] <= matmult_in_a128;
    a[129] <= matmult_in_a129;
    a[130] <= matmult_in_a130;
    a[131] <= matmult_in_a131;
    a[132] <= matmult_in_a132;
    a[133] <= matmult_in_a133;
    a[134] <= matmult_in_a134;
    a[135] <= matmult_in_a135;
    a[136] <= matmult_in_a136;
    a[137] <= matmult_in_a137;
    a[138] <= matmult_in_a138;
    a[139] <= matmult_in_a139;
    a[140] <= matmult_in_a140;
    a[141] <= matmult_in_a141;
    a[142] <= matmult_in_a142;
    a[143] <= matmult_in_a143;
    a[144] <= matmult_in_a144;
    a[145] <= matmult_in_a145;
    a[146] <= matmult_in_a146;
    a[147] <= matmult_in_a147;
    a[148] <= matmult_in_a148;
    a[149] <= matmult_in_a149;
    a[150] <= matmult_in_a150;
    a[151] <= matmult_in_a151;
    a[152] <= matmult_in_a152;
    a[153] <= matmult_in_a153;
    a[154] <= matmult_in_a154;
    a[155] <= matmult_in_a155;
    a[156] <= matmult_in_a156;
    a[157] <= matmult_in_a157;
    a[158] <= matmult_in_a158;
    a[159] <= matmult_in_a159;
    a[160] <= matmult_in_a160;
    a[161] <= matmult_in_a161;
    a[162] <= matmult_in_a162;
    a[163] <= matmult_in_a163;
    a[164] <= matmult_in_a164;
    a[165] <= matmult_in_a165;
    a[166] <= matmult_in_a166;
    a[167] <= matmult_in_a167;
    a[168] <= matmult_in_a168;
    a[169] <= matmult_in_a169;
    a[170] <= matmult_in_a170;
    a[171] <= matmult_in_a171;
    a[172] <= matmult_in_a172;
    a[173] <= matmult_in_a173;
    a[174] <= matmult_in_a174;
    a[175] <= matmult_in_a175;
    a[176] <= matmult_in_a176;
    a[177] <= matmult_in_a177;
    a[178] <= matmult_in_a178;
    a[179] <= matmult_in_a179;
    a[180] <= matmult_in_a180;
    a[181] <= matmult_in_a181;
    a[182] <= matmult_in_a182;
    a[183] <= matmult_in_a183;
    a[184] <= matmult_in_a184;
    a[185] <= matmult_in_a185;
    a[186] <= matmult_in_a186;
    a[187] <= matmult_in_a187;
    a[188] <= matmult_in_a188;
    a[189] <= matmult_in_a189;
    a[190] <= matmult_in_a190;
    a[191] <= matmult_in_a191;
    a[192] <= matmult_in_a192;
    a[193] <= matmult_in_a193;
    a[194] <= matmult_in_a194;
    a[195] <= matmult_in_a195;
    a[196] <= matmult_in_a196;
    a[197] <= matmult_in_a197;
    a[198] <= matmult_in_a198;
    a[199] <= matmult_in_a199;
    a[200] <= matmult_in_a200;
    a[201] <= matmult_in_a201;
    a[202] <= matmult_in_a202;
    a[203] <= matmult_in_a203;
    a[204] <= matmult_in_a204;
    a[205] <= matmult_in_a205;
    a[206] <= matmult_in_a206;
    a[207] <= matmult_in_a207;
    a[208] <= matmult_in_a208;
    a[209] <= matmult_in_a209;
    a[210] <= matmult_in_a210;
    a[211] <= matmult_in_a211;
    a[212] <= matmult_in_a212;
    a[213] <= matmult_in_a213;
    a[214] <= matmult_in_a214;
    a[215] <= matmult_in_a215;
    a[216] <= matmult_in_a216;
    a[217] <= matmult_in_a217;
    a[218] <= matmult_in_a218;
    a[219] <= matmult_in_a219;
    a[220] <= matmult_in_a220;
    a[221] <= matmult_in_a221;
    a[222] <= matmult_in_a222;
    a[223] <= matmult_in_a223;
    a[224] <= matmult_in_a224;
    a[225] <= matmult_in_a225;
    a[226] <= matmult_in_a226;
    a[227] <= matmult_in_a227;
    a[228] <= matmult_in_a228;
    a[229] <= matmult_in_a229;
    a[230] <= matmult_in_a230;
    a[231] <= matmult_in_a231;
    a[232] <= matmult_in_a232;
    a[233] <= matmult_in_a233;
    a[234] <= matmult_in_a234;
    a[235] <= matmult_in_a235;
    a[236] <= matmult_in_a236;
    a[237] <= matmult_in_a237;
    a[238] <= matmult_in_a238;
    a[239] <= matmult_in_a239;
    a[240] <= matmult_in_a240;
    a[241] <= matmult_in_a241;
    a[242] <= matmult_in_a242;
    a[243] <= matmult_in_a243;
    a[244] <= matmult_in_a244;
    a[245] <= matmult_in_a245;
    a[246] <= matmult_in_a246;
    a[247] <= matmult_in_a247;
    a[248] <= matmult_in_a248;
    a[249] <= matmult_in_a249;
    a[250] <= matmult_in_a250;
    a[251] <= matmult_in_a251;
    a[252] <= matmult_in_a252;
    a[253] <= matmult_in_a253;
    a[254] <= matmult_in_a254;
    a[255] <= matmult_in_a255;
    a[256] <= matmult_in_a256;
    a[257] <= matmult_in_a257;
    a[258] <= matmult_in_a258;
    a[259] <= matmult_in_a259;
    a[260] <= matmult_in_a260;
    a[261] <= matmult_in_a261;
    a[262] <= matmult_in_a262;
    a[263] <= matmult_in_a263;
    a[264] <= matmult_in_a264;
    a[265] <= matmult_in_a265;
    a[266] <= matmult_in_a266;
    a[267] <= matmult_in_a267;
    a[268] <= matmult_in_a268;
    a[269] <= matmult_in_a269;
    a[270] <= matmult_in_a270;
    a[271] <= matmult_in_a271;
    a[272] <= matmult_in_a272;
    a[273] <= matmult_in_a273;
    a[274] <= matmult_in_a274;
    a[275] <= matmult_in_a275;
    a[276] <= matmult_in_a276;
    a[277] <= matmult_in_a277;
    a[278] <= matmult_in_a278;
    a[279] <= matmult_in_a279;
    b[0] <= matmult_in_b0;
    b[1] <= matmult_in_b1;
    b[2] <= matmult_in_b2;
    b[3] <= matmult_in_b3;
    b[4] <= matmult_in_b4;
    b[5] <= matmult_in_b5;
    b[6] <= matmult_in_b6;
    b[7] <= matmult_in_b7;
    b[8] <= matmult_in_b8;
    b[9] <= matmult_in_b9;
    b[10] <= matmult_in_b10;
    b[11] <= matmult_in_b11;
    b[12] <= matmult_in_b12;
    b[13] <= matmult_in_b13;
    b[14] <= matmult_in_b14;
    b[15] <= matmult_in_b15;
    b[16] <= matmult_in_b16;
    b[17] <= matmult_in_b17;
    b[18] <= matmult_in_b18;
    b[19] <= matmult_in_b19;
    b[20] <= matmult_in_b20;
    b[21] <= matmult_in_b21;
    b[22] <= matmult_in_b22;
    b[23] <= matmult_in_b23;
    b[24] <= matmult_in_b24;
    b[25] <= matmult_in_b25;
    b[26] <= matmult_in_b26;
    b[27] <= matmult_in_b27;
    b[28] <= matmult_in_b28;
    b[29] <= matmult_in_b29;
    b[30] <= matmult_in_b30;
    b[31] <= matmult_in_b31;
    b[32] <= matmult_in_b32;
    b[33] <= matmult_in_b33;
    b[34] <= matmult_in_b34;
    b[35] <= matmult_in_b35;
    b[36] <= matmult_in_b36;
    b[37] <= matmult_in_b37;
    b[38] <= matmult_in_b38;
    b[39] <= matmult_in_b39;
    b[40] <= matmult_in_b40;
    b[41] <= matmult_in_b41;
    b[42] <= matmult_in_b42;
    b[43] <= matmult_in_b43;
    b[44] <= matmult_in_b44;
    b[45] <= matmult_in_b45;
    b[46] <= matmult_in_b46;
    b[47] <= matmult_in_b47;
    b[48] <= matmult_in_b48;
    b[49] <= matmult_in_b49;
    b[50] <= matmult_in_b50;
    b[51] <= matmult_in_b51;
    b[52] <= matmult_in_b52;
    b[53] <= matmult_in_b53;
    b[54] <= matmult_in_b54;
    b[55] <= matmult_in_b55;
    b[56] <= matmult_in_b56;
    b[57] <= matmult_in_b57;
    b[58] <= matmult_in_b58;
    b[59] <= matmult_in_b59;
    b[60] <= matmult_in_b60;
    b[61] <= matmult_in_b61;
    b[62] <= matmult_in_b62;
    b[63] <= matmult_in_b63;
    b[64] <= matmult_in_b64;
    b[65] <= matmult_in_b65;
    b[66] <= matmult_in_b66;
    b[67] <= matmult_in_b67;
    b[68] <= matmult_in_b68;
    b[69] <= matmult_in_b69;
    b[70] <= matmult_in_b70;
    b[71] <= matmult_in_b71;
    b[72] <= matmult_in_b72;
    b[73] <= matmult_in_b73;
    b[74] <= matmult_in_b74;
    b[75] <= matmult_in_b75;
    b[76] <= matmult_in_b76;
    b[77] <= matmult_in_b77;
    b[78] <= matmult_in_b78;
    b[79] <= matmult_in_b79;
    b[80] <= matmult_in_b80;
    b[81] <= matmult_in_b81;
    b[82] <= matmult_in_b82;
    b[83] <= matmult_in_b83;
    b[84] <= matmult_in_b84;
    b[85] <= matmult_in_b85;
    b[86] <= matmult_in_b86;
    b[87] <= matmult_in_b87;
    b[88] <= matmult_in_b88;
    b[89] <= matmult_in_b89;
    b[90] <= matmult_in_b90;
    b[91] <= matmult_in_b91;
    b[92] <= matmult_in_b92;
    b[93] <= matmult_in_b93;
    b[94] <= matmult_in_b94;
    b[95] <= matmult_in_b95;
    b[96] <= matmult_in_b96;
    b[97] <= matmult_in_b97;
    b[98] <= matmult_in_b98;
    b[99] <= matmult_in_b99;
    b[100] <= matmult_in_b100;
    b[101] <= matmult_in_b101;
    b[102] <= matmult_in_b102;
    b[103] <= matmult_in_b103;
    b[104] <= matmult_in_b104;
    b[105] <= matmult_in_b105;
    b[106] <= matmult_in_b106;
    b[107] <= matmult_in_b107;
    b[108] <= matmult_in_b108;
    b[109] <= matmult_in_b109;
    b[110] <= matmult_in_b110;
    b[111] <= matmult_in_b111;
    b[112] <= matmult_in_b112;
    b[113] <= matmult_in_b113;
    b[114] <= matmult_in_b114;
    b[115] <= matmult_in_b115;
    b[116] <= matmult_in_b116;
    b[117] <= matmult_in_b117;
    b[118] <= matmult_in_b118;
    b[119] <= matmult_in_b119;
    b[120] <= matmult_in_b120;
    b[121] <= matmult_in_b121;
    b[122] <= matmult_in_b122;
    b[123] <= matmult_in_b123;
    b[124] <= matmult_in_b124;
    b[125] <= matmult_in_b125;
    b[126] <= matmult_in_b126;
    b[127] <= matmult_in_b127;
    b[128] <= matmult_in_b128;
    b[129] <= matmult_in_b129;
    b[130] <= matmult_in_b130;
    b[131] <= matmult_in_b131;
    b[132] <= matmult_in_b132;
    b[133] <= matmult_in_b133;
    b[134] <= matmult_in_b134;
    b[135] <= matmult_in_b135;
    b[136] <= matmult_in_b136;
    b[137] <= matmult_in_b137;
    b[138] <= matmult_in_b138;
    b[139] <= matmult_in_b139;
    b[140] <= matmult_in_b140;
    b[141] <= matmult_in_b141;
    b[142] <= matmult_in_b142;
    b[143] <= matmult_in_b143;
    b[144] <= matmult_in_b144;
    b[145] <= matmult_in_b145;
    b[146] <= matmult_in_b146;
    b[147] <= matmult_in_b147;
    b[148] <= matmult_in_b148;
    b[149] <= matmult_in_b149;
    b[150] <= matmult_in_b150;
    b[151] <= matmult_in_b151;
    b[152] <= matmult_in_b152;
    b[153] <= matmult_in_b153;
    b[154] <= matmult_in_b154;
    b[155] <= matmult_in_b155;
    b[156] <= matmult_in_b156;
    b[157] <= matmult_in_b157;
    b[158] <= matmult_in_b158;
    b[159] <= matmult_in_b159;
    b[160] <= matmult_in_b160;
    b[161] <= matmult_in_b161;
    b[162] <= matmult_in_b162;
    b[163] <= matmult_in_b163;
    b[164] <= matmult_in_b164;
    b[165] <= matmult_in_b165;
    b[166] <= matmult_in_b166;
    b[167] <= matmult_in_b167;
    b[168] <= matmult_in_b168;
    b[169] <= matmult_in_b169;
    b[170] <= matmult_in_b170;
    b[171] <= matmult_in_b171;
    b[172] <= matmult_in_b172;
    b[173] <= matmult_in_b173;
    b[174] <= matmult_in_b174;
    b[175] <= matmult_in_b175;
    b[176] <= matmult_in_b176;
    b[177] <= matmult_in_b177;
    b[178] <= matmult_in_b178;
    b[179] <= matmult_in_b179;
    b[180] <= matmult_in_b180;
    b[181] <= matmult_in_b181;
    b[182] <= matmult_in_b182;
    b[183] <= matmult_in_b183;
    b[184] <= matmult_in_b184;
    b[185] <= matmult_in_b185;
    b[186] <= matmult_in_b186;
    b[187] <= matmult_in_b187;
    b[188] <= matmult_in_b188;
    b[189] <= matmult_in_b189;
    b[190] <= matmult_in_b190;
    b[191] <= matmult_in_b191;
    b[192] <= matmult_in_b192;
    b[193] <= matmult_in_b193;
    b[194] <= matmult_in_b194;
    b[195] <= matmult_in_b195;
    b[196] <= matmult_in_b196;
    b[197] <= matmult_in_b197;
    b[198] <= matmult_in_b198;
    b[199] <= matmult_in_b199;
    b[200] <= matmult_in_b200;
    b[201] <= matmult_in_b201;
    b[202] <= matmult_in_b202;
    b[203] <= matmult_in_b203;
    b[204] <= matmult_in_b204;
    b[205] <= matmult_in_b205;
    b[206] <= matmult_in_b206;
    b[207] <= matmult_in_b207;
    b[208] <= matmult_in_b208;
    b[209] <= matmult_in_b209;
    b[210] <= matmult_in_b210;
    b[211] <= matmult_in_b211;
    b[212] <= matmult_in_b212;
    b[213] <= matmult_in_b213;
    b[214] <= matmult_in_b214;
    b[215] <= matmult_in_b215;
    b[216] <= matmult_in_b216;
    b[217] <= matmult_in_b217;
    b[218] <= matmult_in_b218;
    b[219] <= matmult_in_b219;
    b[220] <= matmult_in_b220;
    b[221] <= matmult_in_b221;
    b[222] <= matmult_in_b222;
    b[223] <= matmult_in_b223;
    b[224] <= matmult_in_b224;
    b[225] <= matmult_in_b225;
    b[226] <= matmult_in_b226;
    b[227] <= matmult_in_b227;
    b[228] <= matmult_in_b228;
    b[229] <= matmult_in_b229;
    b[230] <= matmult_in_b230;
    b[231] <= matmult_in_b231;
    b[232] <= matmult_in_b232;
    b[233] <= matmult_in_b233;
    b[234] <= matmult_in_b234;
    b[235] <= matmult_in_b235;
    b[236] <= matmult_in_b236;
    b[237] <= matmult_in_b237;
    b[238] <= matmult_in_b238;
    b[239] <= matmult_in_b239;
    b[240] <= matmult_in_b240;
    b[241] <= matmult_in_b241;
    b[242] <= matmult_in_b242;
    b[243] <= matmult_in_b243;
    b[244] <= matmult_in_b244;
    b[245] <= matmult_in_b245;
    b[246] <= matmult_in_b246;
    b[247] <= matmult_in_b247;
    b[248] <= matmult_in_b248;
    b[249] <= matmult_in_b249;
    b[250] <= matmult_in_b250;
    b[251] <= matmult_in_b251;
    b[252] <= matmult_in_b252;
    b[253] <= matmult_in_b253;
    b[254] <= matmult_in_b254;
    b[255] <= matmult_in_b255;
    b[256] <= matmult_in_b256;
    b[257] <= matmult_in_b257;
    b[258] <= matmult_in_b258;
    b[259] <= matmult_in_b259;
    b[260] <= matmult_in_b260;
    b[261] <= matmult_in_b261;
    b[262] <= matmult_in_b262;
    b[263] <= matmult_in_b263;
    b[264] <= matmult_in_b264;
    b[265] <= matmult_in_b265;
    b[266] <= matmult_in_b266;
    b[267] <= matmult_in_b267;
    b[268] <= matmult_in_b268;
    b[269] <= matmult_in_b269;
    b[270] <= matmult_in_b270;
    b[271] <= matmult_in_b271;
    b[272] <= matmult_in_b272;
    b[273] <= matmult_in_b273;
    b[274] <= matmult_in_b274;
    b[275] <= matmult_in_b275;
    b[276] <= matmult_in_b276;
    b[277] <= matmult_in_b277;
    b[278] <= matmult_in_b278;
    b[279] <= matmult_in_b279;
end

                end
                fin: begin
                    matmult_valid <= 1;
                end
                calc: begin
                    c[0] <= a[0] * b[0] + a[1] * b[14] + a[2] * b[28] + a[3] * b[42] + a[4] * b[56] + a[5] * b[70] + a[6] * b[84] + a[7] * b[98] + a[8] * b[112] + a[9] * b[126] + a[10] * b[140] + a[11] * b[154] + a[12] * b[168] + a[13] * b[182];
                    c[1] <= a[0] * b[1] + a[1] * b[15] + a[2] * b[29] + a[3] * b[43] + a[4] * b[57] + a[5] * b[71] + a[6] * b[85] + a[7] * b[99] + a[8] * b[113] + a[9] * b[127] + a[10] * b[141] + a[11] * b[155] + a[12] * b[169] + a[13] * b[183];
                    c[2] <= a[0] * b[2] + a[1] * b[16] + a[2] * b[30] + a[3] * b[44] + a[4] * b[58] + a[5] * b[72] + a[6] * b[86] + a[7] * b[100] + a[8] * b[114] + a[9] * b[128] + a[10] * b[142] + a[11] * b[156] + a[12] * b[170] + a[13] * b[184];
                    c[3] <= a[0] * b[3] + a[1] * b[17] + a[2] * b[31] + a[3] * b[45] + a[4] * b[59] + a[5] * b[73] + a[6] * b[87] + a[7] * b[101] + a[8] * b[115] + a[9] * b[129] + a[10] * b[143] + a[11] * b[157] + a[12] * b[171] + a[13] * b[185];
                    c[4] <= a[0] * b[4] + a[1] * b[18] + a[2] * b[32] + a[3] * b[46] + a[4] * b[60] + a[5] * b[74] + a[6] * b[88] + a[7] * b[102] + a[8] * b[116] + a[9] * b[130] + a[10] * b[144] + a[11] * b[158] + a[12] * b[172] + a[13] * b[186];
                    c[5] <= a[0] * b[5] + a[1] * b[19] + a[2] * b[33] + a[3] * b[47] + a[4] * b[61] + a[5] * b[75] + a[6] * b[89] + a[7] * b[103] + a[8] * b[117] + a[9] * b[131] + a[10] * b[145] + a[11] * b[159] + a[12] * b[173] + a[13] * b[187];
                    c[6] <= a[0] * b[6] + a[1] * b[20] + a[2] * b[34] + a[3] * b[48] + a[4] * b[62] + a[5] * b[76] + a[6] * b[90] + a[7] * b[104] + a[8] * b[118] + a[9] * b[132] + a[10] * b[146] + a[11] * b[160] + a[12] * b[174] + a[13] * b[188];
                    c[7] <= a[0] * b[7] + a[1] * b[21] + a[2] * b[35] + a[3] * b[49] + a[4] * b[63] + a[5] * b[77] + a[6] * b[91] + a[7] * b[105] + a[8] * b[119] + a[9] * b[133] + a[10] * b[147] + a[11] * b[161] + a[12] * b[175] + a[13] * b[189];
                    c[8] <= a[0] * b[8] + a[1] * b[22] + a[2] * b[36] + a[3] * b[50] + a[4] * b[64] + a[5] * b[78] + a[6] * b[92] + a[7] * b[106] + a[8] * b[120] + a[9] * b[134] + a[10] * b[148] + a[11] * b[162] + a[12] * b[176] + a[13] * b[190];
                    c[9] <= a[0] * b[9] + a[1] * b[23] + a[2] * b[37] + a[3] * b[51] + a[4] * b[65] + a[5] * b[79] + a[6] * b[93] + a[7] * b[107] + a[8] * b[121] + a[9] * b[135] + a[10] * b[149] + a[11] * b[163] + a[12] * b[177] + a[13] * b[191];
                    c[10] <= a[0] * b[10] + a[1] * b[24] + a[2] * b[38] + a[3] * b[52] + a[4] * b[66] + a[5] * b[80] + a[6] * b[94] + a[7] * b[108] + a[8] * b[122] + a[9] * b[136] + a[10] * b[150] + a[11] * b[164] + a[12] * b[178] + a[13] * b[192];
                    c[11] <= a[0] * b[11] + a[1] * b[25] + a[2] * b[39] + a[3] * b[53] + a[4] * b[67] + a[5] * b[81] + a[6] * b[95] + a[7] * b[109] + a[8] * b[123] + a[9] * b[137] + a[10] * b[151] + a[11] * b[165] + a[12] * b[179] + a[13] * b[193];
                    c[12] <= a[0] * b[12] + a[1] * b[26] + a[2] * b[40] + a[3] * b[54] + a[4] * b[68] + a[5] * b[82] + a[6] * b[96] + a[7] * b[110] + a[8] * b[124] + a[9] * b[138] + a[10] * b[152] + a[11] * b[166] + a[12] * b[180] + a[13] * b[194];
                    c[13] <= a[0] * b[13] + a[1] * b[27] + a[2] * b[41] + a[3] * b[55] + a[4] * b[69] + a[5] * b[83] + a[6] * b[97] + a[7] * b[111] + a[8] * b[125] + a[9] * b[139] + a[10] * b[153] + a[11] * b[167] + a[12] * b[181] + a[13] * b[195];
                    c[14] <= a[14] * b[0] + a[15] * b[14] + a[16] * b[28] + a[17] * b[42] + a[18] * b[56] + a[19] * b[70] + a[20] * b[84] + a[21] * b[98] + a[22] * b[112] + a[23] * b[126] + a[24] * b[140] + a[25] * b[154] + a[26] * b[168] + a[27] * b[182];
                    c[15] <= a[14] * b[1] + a[15] * b[15] + a[16] * b[29] + a[17] * b[43] + a[18] * b[57] + a[19] * b[71] + a[20] * b[85] + a[21] * b[99] + a[22] * b[113] + a[23] * b[127] + a[24] * b[141] + a[25] * b[155] + a[26] * b[169] + a[27] * b[183];
                    c[16] <= a[14] * b[2] + a[15] * b[16] + a[16] * b[30] + a[17] * b[44] + a[18] * b[58] + a[19] * b[72] + a[20] * b[86] + a[21] * b[100] + a[22] * b[114] + a[23] * b[128] + a[24] * b[142] + a[25] * b[156] + a[26] * b[170] + a[27] * b[184];
                    c[17] <= a[14] * b[3] + a[15] * b[17] + a[16] * b[31] + a[17] * b[45] + a[18] * b[59] + a[19] * b[73] + a[20] * b[87] + a[21] * b[101] + a[22] * b[115] + a[23] * b[129] + a[24] * b[143] + a[25] * b[157] + a[26] * b[171] + a[27] * b[185];
                    c[18] <= a[14] * b[4] + a[15] * b[18] + a[16] * b[32] + a[17] * b[46] + a[18] * b[60] + a[19] * b[74] + a[20] * b[88] + a[21] * b[102] + a[22] * b[116] + a[23] * b[130] + a[24] * b[144] + a[25] * b[158] + a[26] * b[172] + a[27] * b[186];
                    c[19] <= a[14] * b[5] + a[15] * b[19] + a[16] * b[33] + a[17] * b[47] + a[18] * b[61] + a[19] * b[75] + a[20] * b[89] + a[21] * b[103] + a[22] * b[117] + a[23] * b[131] + a[24] * b[145] + a[25] * b[159] + a[26] * b[173] + a[27] * b[187];
                    c[20] <= a[14] * b[6] + a[15] * b[20] + a[16] * b[34] + a[17] * b[48] + a[18] * b[62] + a[19] * b[76] + a[20] * b[90] + a[21] * b[104] + a[22] * b[118] + a[23] * b[132] + a[24] * b[146] + a[25] * b[160] + a[26] * b[174] + a[27] * b[188];
                    c[21] <= a[14] * b[7] + a[15] * b[21] + a[16] * b[35] + a[17] * b[49] + a[18] * b[63] + a[19] * b[77] + a[20] * b[91] + a[21] * b[105] + a[22] * b[119] + a[23] * b[133] + a[24] * b[147] + a[25] * b[161] + a[26] * b[175] + a[27] * b[189];
                    c[22] <= a[14] * b[8] + a[15] * b[22] + a[16] * b[36] + a[17] * b[50] + a[18] * b[64] + a[19] * b[78] + a[20] * b[92] + a[21] * b[106] + a[22] * b[120] + a[23] * b[134] + a[24] * b[148] + a[25] * b[162] + a[26] * b[176] + a[27] * b[190];
                    c[23] <= a[14] * b[9] + a[15] * b[23] + a[16] * b[37] + a[17] * b[51] + a[18] * b[65] + a[19] * b[79] + a[20] * b[93] + a[21] * b[107] + a[22] * b[121] + a[23] * b[135] + a[24] * b[149] + a[25] * b[163] + a[26] * b[177] + a[27] * b[191];
                    c[24] <= a[14] * b[10] + a[15] * b[24] + a[16] * b[38] + a[17] * b[52] + a[18] * b[66] + a[19] * b[80] + a[20] * b[94] + a[21] * b[108] + a[22] * b[122] + a[23] * b[136] + a[24] * b[150] + a[25] * b[164] + a[26] * b[178] + a[27] * b[192];
                    c[25] <= a[14] * b[11] + a[15] * b[25] + a[16] * b[39] + a[17] * b[53] + a[18] * b[67] + a[19] * b[81] + a[20] * b[95] + a[21] * b[109] + a[22] * b[123] + a[23] * b[137] + a[24] * b[151] + a[25] * b[165] + a[26] * b[179] + a[27] * b[193];
                    c[26] <= a[14] * b[12] + a[15] * b[26] + a[16] * b[40] + a[17] * b[54] + a[18] * b[68] + a[19] * b[82] + a[20] * b[96] + a[21] * b[110] + a[22] * b[124] + a[23] * b[138] + a[24] * b[152] + a[25] * b[166] + a[26] * b[180] + a[27] * b[194];
                    c[27] <= a[14] * b[13] + a[15] * b[27] + a[16] * b[41] + a[17] * b[55] + a[18] * b[69] + a[19] * b[83] + a[20] * b[97] + a[21] * b[111] + a[22] * b[125] + a[23] * b[139] + a[24] * b[153] + a[25] * b[167] + a[26] * b[181] + a[27] * b[195];
                    c[28] <= a[28] * b[0] + a[29] * b[14] + a[30] * b[28] + a[31] * b[42] + a[32] * b[56] + a[33] * b[70] + a[34] * b[84] + a[35] * b[98] + a[36] * b[112] + a[37] * b[126] + a[38] * b[140] + a[39] * b[154] + a[40] * b[168] + a[41] * b[182];
                    c[29] <= a[28] * b[1] + a[29] * b[15] + a[30] * b[29] + a[31] * b[43] + a[32] * b[57] + a[33] * b[71] + a[34] * b[85] + a[35] * b[99] + a[36] * b[113] + a[37] * b[127] + a[38] * b[141] + a[39] * b[155] + a[40] * b[169] + a[41] * b[183];
                    c[30] <= a[28] * b[2] + a[29] * b[16] + a[30] * b[30] + a[31] * b[44] + a[32] * b[58] + a[33] * b[72] + a[34] * b[86] + a[35] * b[100] + a[36] * b[114] + a[37] * b[128] + a[38] * b[142] + a[39] * b[156] + a[40] * b[170] + a[41] * b[184];
                    c[31] <= a[28] * b[3] + a[29] * b[17] + a[30] * b[31] + a[31] * b[45] + a[32] * b[59] + a[33] * b[73] + a[34] * b[87] + a[35] * b[101] + a[36] * b[115] + a[37] * b[129] + a[38] * b[143] + a[39] * b[157] + a[40] * b[171] + a[41] * b[185];
                    c[32] <= a[28] * b[4] + a[29] * b[18] + a[30] * b[32] + a[31] * b[46] + a[32] * b[60] + a[33] * b[74] + a[34] * b[88] + a[35] * b[102] + a[36] * b[116] + a[37] * b[130] + a[38] * b[144] + a[39] * b[158] + a[40] * b[172] + a[41] * b[186];
                    c[33] <= a[28] * b[5] + a[29] * b[19] + a[30] * b[33] + a[31] * b[47] + a[32] * b[61] + a[33] * b[75] + a[34] * b[89] + a[35] * b[103] + a[36] * b[117] + a[37] * b[131] + a[38] * b[145] + a[39] * b[159] + a[40] * b[173] + a[41] * b[187];
                    c[34] <= a[28] * b[6] + a[29] * b[20] + a[30] * b[34] + a[31] * b[48] + a[32] * b[62] + a[33] * b[76] + a[34] * b[90] + a[35] * b[104] + a[36] * b[118] + a[37] * b[132] + a[38] * b[146] + a[39] * b[160] + a[40] * b[174] + a[41] * b[188];
                    c[35] <= a[28] * b[7] + a[29] * b[21] + a[30] * b[35] + a[31] * b[49] + a[32] * b[63] + a[33] * b[77] + a[34] * b[91] + a[35] * b[105] + a[36] * b[119] + a[37] * b[133] + a[38] * b[147] + a[39] * b[161] + a[40] * b[175] + a[41] * b[189];
                    c[36] <= a[28] * b[8] + a[29] * b[22] + a[30] * b[36] + a[31] * b[50] + a[32] * b[64] + a[33] * b[78] + a[34] * b[92] + a[35] * b[106] + a[36] * b[120] + a[37] * b[134] + a[38] * b[148] + a[39] * b[162] + a[40] * b[176] + a[41] * b[190];
                    c[37] <= a[28] * b[9] + a[29] * b[23] + a[30] * b[37] + a[31] * b[51] + a[32] * b[65] + a[33] * b[79] + a[34] * b[93] + a[35] * b[107] + a[36] * b[121] + a[37] * b[135] + a[38] * b[149] + a[39] * b[163] + a[40] * b[177] + a[41] * b[191];
                    c[38] <= a[28] * b[10] + a[29] * b[24] + a[30] * b[38] + a[31] * b[52] + a[32] * b[66] + a[33] * b[80] + a[34] * b[94] + a[35] * b[108] + a[36] * b[122] + a[37] * b[136] + a[38] * b[150] + a[39] * b[164] + a[40] * b[178] + a[41] * b[192];
                    c[39] <= a[28] * b[11] + a[29] * b[25] + a[30] * b[39] + a[31] * b[53] + a[32] * b[67] + a[33] * b[81] + a[34] * b[95] + a[35] * b[109] + a[36] * b[123] + a[37] * b[137] + a[38] * b[151] + a[39] * b[165] + a[40] * b[179] + a[41] * b[193];
                    c[40] <= a[28] * b[12] + a[29] * b[26] + a[30] * b[40] + a[31] * b[54] + a[32] * b[68] + a[33] * b[82] + a[34] * b[96] + a[35] * b[110] + a[36] * b[124] + a[37] * b[138] + a[38] * b[152] + a[39] * b[166] + a[40] * b[180] + a[41] * b[194];
                    c[41] <= a[28] * b[13] + a[29] * b[27] + a[30] * b[41] + a[31] * b[55] + a[32] * b[69] + a[33] * b[83] + a[34] * b[97] + a[35] * b[111] + a[36] * b[125] + a[37] * b[139] + a[38] * b[153] + a[39] * b[167] + a[40] * b[181] + a[41] * b[195];
                    c[42] <= a[42] * b[0] + a[43] * b[14] + a[44] * b[28] + a[45] * b[42] + a[46] * b[56] + a[47] * b[70] + a[48] * b[84] + a[49] * b[98] + a[50] * b[112] + a[51] * b[126] + a[52] * b[140] + a[53] * b[154] + a[54] * b[168] + a[55] * b[182];
                    c[43] <= a[42] * b[1] + a[43] * b[15] + a[44] * b[29] + a[45] * b[43] + a[46] * b[57] + a[47] * b[71] + a[48] * b[85] + a[49] * b[99] + a[50] * b[113] + a[51] * b[127] + a[52] * b[141] + a[53] * b[155] + a[54] * b[169] + a[55] * b[183];
                    c[44] <= a[42] * b[2] + a[43] * b[16] + a[44] * b[30] + a[45] * b[44] + a[46] * b[58] + a[47] * b[72] + a[48] * b[86] + a[49] * b[100] + a[50] * b[114] + a[51] * b[128] + a[52] * b[142] + a[53] * b[156] + a[54] * b[170] + a[55] * b[184];
                    c[45] <= a[42] * b[3] + a[43] * b[17] + a[44] * b[31] + a[45] * b[45] + a[46] * b[59] + a[47] * b[73] + a[48] * b[87] + a[49] * b[101] + a[50] * b[115] + a[51] * b[129] + a[52] * b[143] + a[53] * b[157] + a[54] * b[171] + a[55] * b[185];
                    c[46] <= a[42] * b[4] + a[43] * b[18] + a[44] * b[32] + a[45] * b[46] + a[46] * b[60] + a[47] * b[74] + a[48] * b[88] + a[49] * b[102] + a[50] * b[116] + a[51] * b[130] + a[52] * b[144] + a[53] * b[158] + a[54] * b[172] + a[55] * b[186];
                    c[47] <= a[42] * b[5] + a[43] * b[19] + a[44] * b[33] + a[45] * b[47] + a[46] * b[61] + a[47] * b[75] + a[48] * b[89] + a[49] * b[103] + a[50] * b[117] + a[51] * b[131] + a[52] * b[145] + a[53] * b[159] + a[54] * b[173] + a[55] * b[187];
                    c[48] <= a[42] * b[6] + a[43] * b[20] + a[44] * b[34] + a[45] * b[48] + a[46] * b[62] + a[47] * b[76] + a[48] * b[90] + a[49] * b[104] + a[50] * b[118] + a[51] * b[132] + a[52] * b[146] + a[53] * b[160] + a[54] * b[174] + a[55] * b[188];
                    c[49] <= a[42] * b[7] + a[43] * b[21] + a[44] * b[35] + a[45] * b[49] + a[46] * b[63] + a[47] * b[77] + a[48] * b[91] + a[49] * b[105] + a[50] * b[119] + a[51] * b[133] + a[52] * b[147] + a[53] * b[161] + a[54] * b[175] + a[55] * b[189];
                    c[50] <= a[42] * b[8] + a[43] * b[22] + a[44] * b[36] + a[45] * b[50] + a[46] * b[64] + a[47] * b[78] + a[48] * b[92] + a[49] * b[106] + a[50] * b[120] + a[51] * b[134] + a[52] * b[148] + a[53] * b[162] + a[54] * b[176] + a[55] * b[190];
                    c[51] <= a[42] * b[9] + a[43] * b[23] + a[44] * b[37] + a[45] * b[51] + a[46] * b[65] + a[47] * b[79] + a[48] * b[93] + a[49] * b[107] + a[50] * b[121] + a[51] * b[135] + a[52] * b[149] + a[53] * b[163] + a[54] * b[177] + a[55] * b[191];
                    c[52] <= a[42] * b[10] + a[43] * b[24] + a[44] * b[38] + a[45] * b[52] + a[46] * b[66] + a[47] * b[80] + a[48] * b[94] + a[49] * b[108] + a[50] * b[122] + a[51] * b[136] + a[52] * b[150] + a[53] * b[164] + a[54] * b[178] + a[55] * b[192];
                    c[53] <= a[42] * b[11] + a[43] * b[25] + a[44] * b[39] + a[45] * b[53] + a[46] * b[67] + a[47] * b[81] + a[48] * b[95] + a[49] * b[109] + a[50] * b[123] + a[51] * b[137] + a[52] * b[151] + a[53] * b[165] + a[54] * b[179] + a[55] * b[193];
                    c[54] <= a[42] * b[12] + a[43] * b[26] + a[44] * b[40] + a[45] * b[54] + a[46] * b[68] + a[47] * b[82] + a[48] * b[96] + a[49] * b[110] + a[50] * b[124] + a[51] * b[138] + a[52] * b[152] + a[53] * b[166] + a[54] * b[180] + a[55] * b[194];
                    c[55] <= a[42] * b[13] + a[43] * b[27] + a[44] * b[41] + a[45] * b[55] + a[46] * b[69] + a[47] * b[83] + a[48] * b[97] + a[49] * b[111] + a[50] * b[125] + a[51] * b[139] + a[52] * b[153] + a[53] * b[167] + a[54] * b[181] + a[55] * b[195];
                    c[56] <= a[56] * b[0] + a[57] * b[14] + a[58] * b[28] + a[59] * b[42] + a[60] * b[56] + a[61] * b[70] + a[62] * b[84] + a[63] * b[98] + a[64] * b[112] + a[65] * b[126] + a[66] * b[140] + a[67] * b[154] + a[68] * b[168] + a[69] * b[182];
                    c[57] <= a[56] * b[1] + a[57] * b[15] + a[58] * b[29] + a[59] * b[43] + a[60] * b[57] + a[61] * b[71] + a[62] * b[85] + a[63] * b[99] + a[64] * b[113] + a[65] * b[127] + a[66] * b[141] + a[67] * b[155] + a[68] * b[169] + a[69] * b[183];
                    c[58] <= a[56] * b[2] + a[57] * b[16] + a[58] * b[30] + a[59] * b[44] + a[60] * b[58] + a[61] * b[72] + a[62] * b[86] + a[63] * b[100] + a[64] * b[114] + a[65] * b[128] + a[66] * b[142] + a[67] * b[156] + a[68] * b[170] + a[69] * b[184];
                    c[59] <= a[56] * b[3] + a[57] * b[17] + a[58] * b[31] + a[59] * b[45] + a[60] * b[59] + a[61] * b[73] + a[62] * b[87] + a[63] * b[101] + a[64] * b[115] + a[65] * b[129] + a[66] * b[143] + a[67] * b[157] + a[68] * b[171] + a[69] * b[185];
                    c[60] <= a[56] * b[4] + a[57] * b[18] + a[58] * b[32] + a[59] * b[46] + a[60] * b[60] + a[61] * b[74] + a[62] * b[88] + a[63] * b[102] + a[64] * b[116] + a[65] * b[130] + a[66] * b[144] + a[67] * b[158] + a[68] * b[172] + a[69] * b[186];
                    c[61] <= a[56] * b[5] + a[57] * b[19] + a[58] * b[33] + a[59] * b[47] + a[60] * b[61] + a[61] * b[75] + a[62] * b[89] + a[63] * b[103] + a[64] * b[117] + a[65] * b[131] + a[66] * b[145] + a[67] * b[159] + a[68] * b[173] + a[69] * b[187];
                    c[62] <= a[56] * b[6] + a[57] * b[20] + a[58] * b[34] + a[59] * b[48] + a[60] * b[62] + a[61] * b[76] + a[62] * b[90] + a[63] * b[104] + a[64] * b[118] + a[65] * b[132] + a[66] * b[146] + a[67] * b[160] + a[68] * b[174] + a[69] * b[188];
                    c[63] <= a[56] * b[7] + a[57] * b[21] + a[58] * b[35] + a[59] * b[49] + a[60] * b[63] + a[61] * b[77] + a[62] * b[91] + a[63] * b[105] + a[64] * b[119] + a[65] * b[133] + a[66] * b[147] + a[67] * b[161] + a[68] * b[175] + a[69] * b[189];
                    c[64] <= a[56] * b[8] + a[57] * b[22] + a[58] * b[36] + a[59] * b[50] + a[60] * b[64] + a[61] * b[78] + a[62] * b[92] + a[63] * b[106] + a[64] * b[120] + a[65] * b[134] + a[66] * b[148] + a[67] * b[162] + a[68] * b[176] + a[69] * b[190];
                    c[65] <= a[56] * b[9] + a[57] * b[23] + a[58] * b[37] + a[59] * b[51] + a[60] * b[65] + a[61] * b[79] + a[62] * b[93] + a[63] * b[107] + a[64] * b[121] + a[65] * b[135] + a[66] * b[149] + a[67] * b[163] + a[68] * b[177] + a[69] * b[191];
                    c[66] <= a[56] * b[10] + a[57] * b[24] + a[58] * b[38] + a[59] * b[52] + a[60] * b[66] + a[61] * b[80] + a[62] * b[94] + a[63] * b[108] + a[64] * b[122] + a[65] * b[136] + a[66] * b[150] + a[67] * b[164] + a[68] * b[178] + a[69] * b[192];
                    c[67] <= a[56] * b[11] + a[57] * b[25] + a[58] * b[39] + a[59] * b[53] + a[60] * b[67] + a[61] * b[81] + a[62] * b[95] + a[63] * b[109] + a[64] * b[123] + a[65] * b[137] + a[66] * b[151] + a[67] * b[165] + a[68] * b[179] + a[69] * b[193];
                    c[68] <= a[56] * b[12] + a[57] * b[26] + a[58] * b[40] + a[59] * b[54] + a[60] * b[68] + a[61] * b[82] + a[62] * b[96] + a[63] * b[110] + a[64] * b[124] + a[65] * b[138] + a[66] * b[152] + a[67] * b[166] + a[68] * b[180] + a[69] * b[194];
                    c[69] <= a[56] * b[13] + a[57] * b[27] + a[58] * b[41] + a[59] * b[55] + a[60] * b[69] + a[61] * b[83] + a[62] * b[97] + a[63] * b[111] + a[64] * b[125] + a[65] * b[139] + a[66] * b[153] + a[67] * b[167] + a[68] * b[181] + a[69] * b[195];
                    c[70] <= a[70] * b[0] + a[71] * b[14] + a[72] * b[28] + a[73] * b[42] + a[74] * b[56] + a[75] * b[70] + a[76] * b[84] + a[77] * b[98] + a[78] * b[112] + a[79] * b[126] + a[80] * b[140] + a[81] * b[154] + a[82] * b[168] + a[83] * b[182];
                    c[71] <= a[70] * b[1] + a[71] * b[15] + a[72] * b[29] + a[73] * b[43] + a[74] * b[57] + a[75] * b[71] + a[76] * b[85] + a[77] * b[99] + a[78] * b[113] + a[79] * b[127] + a[80] * b[141] + a[81] * b[155] + a[82] * b[169] + a[83] * b[183];
                    c[72] <= a[70] * b[2] + a[71] * b[16] + a[72] * b[30] + a[73] * b[44] + a[74] * b[58] + a[75] * b[72] + a[76] * b[86] + a[77] * b[100] + a[78] * b[114] + a[79] * b[128] + a[80] * b[142] + a[81] * b[156] + a[82] * b[170] + a[83] * b[184];
                    c[73] <= a[70] * b[3] + a[71] * b[17] + a[72] * b[31] + a[73] * b[45] + a[74] * b[59] + a[75] * b[73] + a[76] * b[87] + a[77] * b[101] + a[78] * b[115] + a[79] * b[129] + a[80] * b[143] + a[81] * b[157] + a[82] * b[171] + a[83] * b[185];
                    c[74] <= a[70] * b[4] + a[71] * b[18] + a[72] * b[32] + a[73] * b[46] + a[74] * b[60] + a[75] * b[74] + a[76] * b[88] + a[77] * b[102] + a[78] * b[116] + a[79] * b[130] + a[80] * b[144] + a[81] * b[158] + a[82] * b[172] + a[83] * b[186];
                    c[75] <= a[70] * b[5] + a[71] * b[19] + a[72] * b[33] + a[73] * b[47] + a[74] * b[61] + a[75] * b[75] + a[76] * b[89] + a[77] * b[103] + a[78] * b[117] + a[79] * b[131] + a[80] * b[145] + a[81] * b[159] + a[82] * b[173] + a[83] * b[187];
                    c[76] <= a[70] * b[6] + a[71] * b[20] + a[72] * b[34] + a[73] * b[48] + a[74] * b[62] + a[75] * b[76] + a[76] * b[90] + a[77] * b[104] + a[78] * b[118] + a[79] * b[132] + a[80] * b[146] + a[81] * b[160] + a[82] * b[174] + a[83] * b[188];
                    c[77] <= a[70] * b[7] + a[71] * b[21] + a[72] * b[35] + a[73] * b[49] + a[74] * b[63] + a[75] * b[77] + a[76] * b[91] + a[77] * b[105] + a[78] * b[119] + a[79] * b[133] + a[80] * b[147] + a[81] * b[161] + a[82] * b[175] + a[83] * b[189];
                    c[78] <= a[70] * b[8] + a[71] * b[22] + a[72] * b[36] + a[73] * b[50] + a[74] * b[64] + a[75] * b[78] + a[76] * b[92] + a[77] * b[106] + a[78] * b[120] + a[79] * b[134] + a[80] * b[148] + a[81] * b[162] + a[82] * b[176] + a[83] * b[190];
                    c[79] <= a[70] * b[9] + a[71] * b[23] + a[72] * b[37] + a[73] * b[51] + a[74] * b[65] + a[75] * b[79] + a[76] * b[93] + a[77] * b[107] + a[78] * b[121] + a[79] * b[135] + a[80] * b[149] + a[81] * b[163] + a[82] * b[177] + a[83] * b[191];
                    c[80] <= a[70] * b[10] + a[71] * b[24] + a[72] * b[38] + a[73] * b[52] + a[74] * b[66] + a[75] * b[80] + a[76] * b[94] + a[77] * b[108] + a[78] * b[122] + a[79] * b[136] + a[80] * b[150] + a[81] * b[164] + a[82] * b[178] + a[83] * b[192];
                    c[81] <= a[70] * b[11] + a[71] * b[25] + a[72] * b[39] + a[73] * b[53] + a[74] * b[67] + a[75] * b[81] + a[76] * b[95] + a[77] * b[109] + a[78] * b[123] + a[79] * b[137] + a[80] * b[151] + a[81] * b[165] + a[82] * b[179] + a[83] * b[193];
                    c[82] <= a[70] * b[12] + a[71] * b[26] + a[72] * b[40] + a[73] * b[54] + a[74] * b[68] + a[75] * b[82] + a[76] * b[96] + a[77] * b[110] + a[78] * b[124] + a[79] * b[138] + a[80] * b[152] + a[81] * b[166] + a[82] * b[180] + a[83] * b[194];
                    c[83] <= a[70] * b[13] + a[71] * b[27] + a[72] * b[41] + a[73] * b[55] + a[74] * b[69] + a[75] * b[83] + a[76] * b[97] + a[77] * b[111] + a[78] * b[125] + a[79] * b[139] + a[80] * b[153] + a[81] * b[167] + a[82] * b[181] + a[83] * b[195];
                    c[84] <= a[84] * b[0] + a[85] * b[14] + a[86] * b[28] + a[87] * b[42] + a[88] * b[56] + a[89] * b[70] + a[90] * b[84] + a[91] * b[98] + a[92] * b[112] + a[93] * b[126] + a[94] * b[140] + a[95] * b[154] + a[96] * b[168] + a[97] * b[182];
                    c[85] <= a[84] * b[1] + a[85] * b[15] + a[86] * b[29] + a[87] * b[43] + a[88] * b[57] + a[89] * b[71] + a[90] * b[85] + a[91] * b[99] + a[92] * b[113] + a[93] * b[127] + a[94] * b[141] + a[95] * b[155] + a[96] * b[169] + a[97] * b[183];
                    c[86] <= a[84] * b[2] + a[85] * b[16] + a[86] * b[30] + a[87] * b[44] + a[88] * b[58] + a[89] * b[72] + a[90] * b[86] + a[91] * b[100] + a[92] * b[114] + a[93] * b[128] + a[94] * b[142] + a[95] * b[156] + a[96] * b[170] + a[97] * b[184];
                    c[87] <= a[84] * b[3] + a[85] * b[17] + a[86] * b[31] + a[87] * b[45] + a[88] * b[59] + a[89] * b[73] + a[90] * b[87] + a[91] * b[101] + a[92] * b[115] + a[93] * b[129] + a[94] * b[143] + a[95] * b[157] + a[96] * b[171] + a[97] * b[185];
                    c[88] <= a[84] * b[4] + a[85] * b[18] + a[86] * b[32] + a[87] * b[46] + a[88] * b[60] + a[89] * b[74] + a[90] * b[88] + a[91] * b[102] + a[92] * b[116] + a[93] * b[130] + a[94] * b[144] + a[95] * b[158] + a[96] * b[172] + a[97] * b[186];
                    c[89] <= a[84] * b[5] + a[85] * b[19] + a[86] * b[33] + a[87] * b[47] + a[88] * b[61] + a[89] * b[75] + a[90] * b[89] + a[91] * b[103] + a[92] * b[117] + a[93] * b[131] + a[94] * b[145] + a[95] * b[159] + a[96] * b[173] + a[97] * b[187];
                    c[90] <= a[84] * b[6] + a[85] * b[20] + a[86] * b[34] + a[87] * b[48] + a[88] * b[62] + a[89] * b[76] + a[90] * b[90] + a[91] * b[104] + a[92] * b[118] + a[93] * b[132] + a[94] * b[146] + a[95] * b[160] + a[96] * b[174] + a[97] * b[188];
                    c[91] <= a[84] * b[7] + a[85] * b[21] + a[86] * b[35] + a[87] * b[49] + a[88] * b[63] + a[89] * b[77] + a[90] * b[91] + a[91] * b[105] + a[92] * b[119] + a[93] * b[133] + a[94] * b[147] + a[95] * b[161] + a[96] * b[175] + a[97] * b[189];
                    c[92] <= a[84] * b[8] + a[85] * b[22] + a[86] * b[36] + a[87] * b[50] + a[88] * b[64] + a[89] * b[78] + a[90] * b[92] + a[91] * b[106] + a[92] * b[120] + a[93] * b[134] + a[94] * b[148] + a[95] * b[162] + a[96] * b[176] + a[97] * b[190];
                    c[93] <= a[84] * b[9] + a[85] * b[23] + a[86] * b[37] + a[87] * b[51] + a[88] * b[65] + a[89] * b[79] + a[90] * b[93] + a[91] * b[107] + a[92] * b[121] + a[93] * b[135] + a[94] * b[149] + a[95] * b[163] + a[96] * b[177] + a[97] * b[191];
                    c[94] <= a[84] * b[10] + a[85] * b[24] + a[86] * b[38] + a[87] * b[52] + a[88] * b[66] + a[89] * b[80] + a[90] * b[94] + a[91] * b[108] + a[92] * b[122] + a[93] * b[136] + a[94] * b[150] + a[95] * b[164] + a[96] * b[178] + a[97] * b[192];
                    c[95] <= a[84] * b[11] + a[85] * b[25] + a[86] * b[39] + a[87] * b[53] + a[88] * b[67] + a[89] * b[81] + a[90] * b[95] + a[91] * b[109] + a[92] * b[123] + a[93] * b[137] + a[94] * b[151] + a[95] * b[165] + a[96] * b[179] + a[97] * b[193];
                    c[96] <= a[84] * b[12] + a[85] * b[26] + a[86] * b[40] + a[87] * b[54] + a[88] * b[68] + a[89] * b[82] + a[90] * b[96] + a[91] * b[110] + a[92] * b[124] + a[93] * b[138] + a[94] * b[152] + a[95] * b[166] + a[96] * b[180] + a[97] * b[194];
                    c[97] <= a[84] * b[13] + a[85] * b[27] + a[86] * b[41] + a[87] * b[55] + a[88] * b[69] + a[89] * b[83] + a[90] * b[97] + a[91] * b[111] + a[92] * b[125] + a[93] * b[139] + a[94] * b[153] + a[95] * b[167] + a[96] * b[181] + a[97] * b[195];
                    c[98] <= a[98] * b[0] + a[99] * b[14] + a[100] * b[28] + a[101] * b[42] + a[102] * b[56] + a[103] * b[70] + a[104] * b[84] + a[105] * b[98] + a[106] * b[112] + a[107] * b[126] + a[108] * b[140] + a[109] * b[154] + a[110] * b[168] + a[111] * b[182];
                    c[99] <= a[98] * b[1] + a[99] * b[15] + a[100] * b[29] + a[101] * b[43] + a[102] * b[57] + a[103] * b[71] + a[104] * b[85] + a[105] * b[99] + a[106] * b[113] + a[107] * b[127] + a[108] * b[141] + a[109] * b[155] + a[110] * b[169] + a[111] * b[183];
                    c[100] <= a[98] * b[2] + a[99] * b[16] + a[100] * b[30] + a[101] * b[44] + a[102] * b[58] + a[103] * b[72] + a[104] * b[86] + a[105] * b[100] + a[106] * b[114] + a[107] * b[128] + a[108] * b[142] + a[109] * b[156] + a[110] * b[170] + a[111] * b[184];
                    c[101] <= a[98] * b[3] + a[99] * b[17] + a[100] * b[31] + a[101] * b[45] + a[102] * b[59] + a[103] * b[73] + a[104] * b[87] + a[105] * b[101] + a[106] * b[115] + a[107] * b[129] + a[108] * b[143] + a[109] * b[157] + a[110] * b[171] + a[111] * b[185];
                    c[102] <= a[98] * b[4] + a[99] * b[18] + a[100] * b[32] + a[101] * b[46] + a[102] * b[60] + a[103] * b[74] + a[104] * b[88] + a[105] * b[102] + a[106] * b[116] + a[107] * b[130] + a[108] * b[144] + a[109] * b[158] + a[110] * b[172] + a[111] * b[186];
                    c[103] <= a[98] * b[5] + a[99] * b[19] + a[100] * b[33] + a[101] * b[47] + a[102] * b[61] + a[103] * b[75] + a[104] * b[89] + a[105] * b[103] + a[106] * b[117] + a[107] * b[131] + a[108] * b[145] + a[109] * b[159] + a[110] * b[173] + a[111] * b[187];
                    c[104] <= a[98] * b[6] + a[99] * b[20] + a[100] * b[34] + a[101] * b[48] + a[102] * b[62] + a[103] * b[76] + a[104] * b[90] + a[105] * b[104] + a[106] * b[118] + a[107] * b[132] + a[108] * b[146] + a[109] * b[160] + a[110] * b[174] + a[111] * b[188];
                    c[105] <= a[98] * b[7] + a[99] * b[21] + a[100] * b[35] + a[101] * b[49] + a[102] * b[63] + a[103] * b[77] + a[104] * b[91] + a[105] * b[105] + a[106] * b[119] + a[107] * b[133] + a[108] * b[147] + a[109] * b[161] + a[110] * b[175] + a[111] * b[189];
                    c[106] <= a[98] * b[8] + a[99] * b[22] + a[100] * b[36] + a[101] * b[50] + a[102] * b[64] + a[103] * b[78] + a[104] * b[92] + a[105] * b[106] + a[106] * b[120] + a[107] * b[134] + a[108] * b[148] + a[109] * b[162] + a[110] * b[176] + a[111] * b[190];
                    c[107] <= a[98] * b[9] + a[99] * b[23] + a[100] * b[37] + a[101] * b[51] + a[102] * b[65] + a[103] * b[79] + a[104] * b[93] + a[105] * b[107] + a[106] * b[121] + a[107] * b[135] + a[108] * b[149] + a[109] * b[163] + a[110] * b[177] + a[111] * b[191];
                    c[108] <= a[98] * b[10] + a[99] * b[24] + a[100] * b[38] + a[101] * b[52] + a[102] * b[66] + a[103] * b[80] + a[104] * b[94] + a[105] * b[108] + a[106] * b[122] + a[107] * b[136] + a[108] * b[150] + a[109] * b[164] + a[110] * b[178] + a[111] * b[192];
                    c[109] <= a[98] * b[11] + a[99] * b[25] + a[100] * b[39] + a[101] * b[53] + a[102] * b[67] + a[103] * b[81] + a[104] * b[95] + a[105] * b[109] + a[106] * b[123] + a[107] * b[137] + a[108] * b[151] + a[109] * b[165] + a[110] * b[179] + a[111] * b[193];
                    c[110] <= a[98] * b[12] + a[99] * b[26] + a[100] * b[40] + a[101] * b[54] + a[102] * b[68] + a[103] * b[82] + a[104] * b[96] + a[105] * b[110] + a[106] * b[124] + a[107] * b[138] + a[108] * b[152] + a[109] * b[166] + a[110] * b[180] + a[111] * b[194];
                    c[111] <= a[98] * b[13] + a[99] * b[27] + a[100] * b[41] + a[101] * b[55] + a[102] * b[69] + a[103] * b[83] + a[104] * b[97] + a[105] * b[111] + a[106] * b[125] + a[107] * b[139] + a[108] * b[153] + a[109] * b[167] + a[110] * b[181] + a[111] * b[195];
                    c[112] <= a[112] * b[0] + a[113] * b[14] + a[114] * b[28] + a[115] * b[42] + a[116] * b[56] + a[117] * b[70] + a[118] * b[84] + a[119] * b[98] + a[120] * b[112] + a[121] * b[126] + a[122] * b[140] + a[123] * b[154] + a[124] * b[168] + a[125] * b[182];
                    c[113] <= a[112] * b[1] + a[113] * b[15] + a[114] * b[29] + a[115] * b[43] + a[116] * b[57] + a[117] * b[71] + a[118] * b[85] + a[119] * b[99] + a[120] * b[113] + a[121] * b[127] + a[122] * b[141] + a[123] * b[155] + a[124] * b[169] + a[125] * b[183];
                    c[114] <= a[112] * b[2] + a[113] * b[16] + a[114] * b[30] + a[115] * b[44] + a[116] * b[58] + a[117] * b[72] + a[118] * b[86] + a[119] * b[100] + a[120] * b[114] + a[121] * b[128] + a[122] * b[142] + a[123] * b[156] + a[124] * b[170] + a[125] * b[184];
                    c[115] <= a[112] * b[3] + a[113] * b[17] + a[114] * b[31] + a[115] * b[45] + a[116] * b[59] + a[117] * b[73] + a[118] * b[87] + a[119] * b[101] + a[120] * b[115] + a[121] * b[129] + a[122] * b[143] + a[123] * b[157] + a[124] * b[171] + a[125] * b[185];
                    c[116] <= a[112] * b[4] + a[113] * b[18] + a[114] * b[32] + a[115] * b[46] + a[116] * b[60] + a[117] * b[74] + a[118] * b[88] + a[119] * b[102] + a[120] * b[116] + a[121] * b[130] + a[122] * b[144] + a[123] * b[158] + a[124] * b[172] + a[125] * b[186];
                    c[117] <= a[112] * b[5] + a[113] * b[19] + a[114] * b[33] + a[115] * b[47] + a[116] * b[61] + a[117] * b[75] + a[118] * b[89] + a[119] * b[103] + a[120] * b[117] + a[121] * b[131] + a[122] * b[145] + a[123] * b[159] + a[124] * b[173] + a[125] * b[187];
                    c[118] <= a[112] * b[6] + a[113] * b[20] + a[114] * b[34] + a[115] * b[48] + a[116] * b[62] + a[117] * b[76] + a[118] * b[90] + a[119] * b[104] + a[120] * b[118] + a[121] * b[132] + a[122] * b[146] + a[123] * b[160] + a[124] * b[174] + a[125] * b[188];
                    c[119] <= a[112] * b[7] + a[113] * b[21] + a[114] * b[35] + a[115] * b[49] + a[116] * b[63] + a[117] * b[77] + a[118] * b[91] + a[119] * b[105] + a[120] * b[119] + a[121] * b[133] + a[122] * b[147] + a[123] * b[161] + a[124] * b[175] + a[125] * b[189];
                    c[120] <= a[112] * b[8] + a[113] * b[22] + a[114] * b[36] + a[115] * b[50] + a[116] * b[64] + a[117] * b[78] + a[118] * b[92] + a[119] * b[106] + a[120] * b[120] + a[121] * b[134] + a[122] * b[148] + a[123] * b[162] + a[124] * b[176] + a[125] * b[190];
                    c[121] <= a[112] * b[9] + a[113] * b[23] + a[114] * b[37] + a[115] * b[51] + a[116] * b[65] + a[117] * b[79] + a[118] * b[93] + a[119] * b[107] + a[120] * b[121] + a[121] * b[135] + a[122] * b[149] + a[123] * b[163] + a[124] * b[177] + a[125] * b[191];
                    c[122] <= a[112] * b[10] + a[113] * b[24] + a[114] * b[38] + a[115] * b[52] + a[116] * b[66] + a[117] * b[80] + a[118] * b[94] + a[119] * b[108] + a[120] * b[122] + a[121] * b[136] + a[122] * b[150] + a[123] * b[164] + a[124] * b[178] + a[125] * b[192];
                    c[123] <= a[112] * b[11] + a[113] * b[25] + a[114] * b[39] + a[115] * b[53] + a[116] * b[67] + a[117] * b[81] + a[118] * b[95] + a[119] * b[109] + a[120] * b[123] + a[121] * b[137] + a[122] * b[151] + a[123] * b[165] + a[124] * b[179] + a[125] * b[193];
                    c[124] <= a[112] * b[12] + a[113] * b[26] + a[114] * b[40] + a[115] * b[54] + a[116] * b[68] + a[117] * b[82] + a[118] * b[96] + a[119] * b[110] + a[120] * b[124] + a[121] * b[138] + a[122] * b[152] + a[123] * b[166] + a[124] * b[180] + a[125] * b[194];
                    c[125] <= a[112] * b[13] + a[113] * b[27] + a[114] * b[41] + a[115] * b[55] + a[116] * b[69] + a[117] * b[83] + a[118] * b[97] + a[119] * b[111] + a[120] * b[125] + a[121] * b[139] + a[122] * b[153] + a[123] * b[167] + a[124] * b[181] + a[125] * b[195];
                    c[126] <= a[126] * b[0] + a[127] * b[14] + a[128] * b[28] + a[129] * b[42] + a[130] * b[56] + a[131] * b[70] + a[132] * b[84] + a[133] * b[98] + a[134] * b[112] + a[135] * b[126] + a[136] * b[140] + a[137] * b[154] + a[138] * b[168] + a[139] * b[182];
                    c[127] <= a[126] * b[1] + a[127] * b[15] + a[128] * b[29] + a[129] * b[43] + a[130] * b[57] + a[131] * b[71] + a[132] * b[85] + a[133] * b[99] + a[134] * b[113] + a[135] * b[127] + a[136] * b[141] + a[137] * b[155] + a[138] * b[169] + a[139] * b[183];
                    c[128] <= a[126] * b[2] + a[127] * b[16] + a[128] * b[30] + a[129] * b[44] + a[130] * b[58] + a[131] * b[72] + a[132] * b[86] + a[133] * b[100] + a[134] * b[114] + a[135] * b[128] + a[136] * b[142] + a[137] * b[156] + a[138] * b[170] + a[139] * b[184];
                    c[129] <= a[126] * b[3] + a[127] * b[17] + a[128] * b[31] + a[129] * b[45] + a[130] * b[59] + a[131] * b[73] + a[132] * b[87] + a[133] * b[101] + a[134] * b[115] + a[135] * b[129] + a[136] * b[143] + a[137] * b[157] + a[138] * b[171] + a[139] * b[185];
                    c[130] <= a[126] * b[4] + a[127] * b[18] + a[128] * b[32] + a[129] * b[46] + a[130] * b[60] + a[131] * b[74] + a[132] * b[88] + a[133] * b[102] + a[134] * b[116] + a[135] * b[130] + a[136] * b[144] + a[137] * b[158] + a[138] * b[172] + a[139] * b[186];
                    c[131] <= a[126] * b[5] + a[127] * b[19] + a[128] * b[33] + a[129] * b[47] + a[130] * b[61] + a[131] * b[75] + a[132] * b[89] + a[133] * b[103] + a[134] * b[117] + a[135] * b[131] + a[136] * b[145] + a[137] * b[159] + a[138] * b[173] + a[139] * b[187];
                    c[132] <= a[126] * b[6] + a[127] * b[20] + a[128] * b[34] + a[129] * b[48] + a[130] * b[62] + a[131] * b[76] + a[132] * b[90] + a[133] * b[104] + a[134] * b[118] + a[135] * b[132] + a[136] * b[146] + a[137] * b[160] + a[138] * b[174] + a[139] * b[188];
                    c[133] <= a[126] * b[7] + a[127] * b[21] + a[128] * b[35] + a[129] * b[49] + a[130] * b[63] + a[131] * b[77] + a[132] * b[91] + a[133] * b[105] + a[134] * b[119] + a[135] * b[133] + a[136] * b[147] + a[137] * b[161] + a[138] * b[175] + a[139] * b[189];
                    c[134] <= a[126] * b[8] + a[127] * b[22] + a[128] * b[36] + a[129] * b[50] + a[130] * b[64] + a[131] * b[78] + a[132] * b[92] + a[133] * b[106] + a[134] * b[120] + a[135] * b[134] + a[136] * b[148] + a[137] * b[162] + a[138] * b[176] + a[139] * b[190];
                    c[135] <= a[126] * b[9] + a[127] * b[23] + a[128] * b[37] + a[129] * b[51] + a[130] * b[65] + a[131] * b[79] + a[132] * b[93] + a[133] * b[107] + a[134] * b[121] + a[135] * b[135] + a[136] * b[149] + a[137] * b[163] + a[138] * b[177] + a[139] * b[191];
                    c[136] <= a[126] * b[10] + a[127] * b[24] + a[128] * b[38] + a[129] * b[52] + a[130] * b[66] + a[131] * b[80] + a[132] * b[94] + a[133] * b[108] + a[134] * b[122] + a[135] * b[136] + a[136] * b[150] + a[137] * b[164] + a[138] * b[178] + a[139] * b[192];
                    c[137] <= a[126] * b[11] + a[127] * b[25] + a[128] * b[39] + a[129] * b[53] + a[130] * b[67] + a[131] * b[81] + a[132] * b[95] + a[133] * b[109] + a[134] * b[123] + a[135] * b[137] + a[136] * b[151] + a[137] * b[165] + a[138] * b[179] + a[139] * b[193];
                    c[138] <= a[126] * b[12] + a[127] * b[26] + a[128] * b[40] + a[129] * b[54] + a[130] * b[68] + a[131] * b[82] + a[132] * b[96] + a[133] * b[110] + a[134] * b[124] + a[135] * b[138] + a[136] * b[152] + a[137] * b[166] + a[138] * b[180] + a[139] * b[194];
                    c[139] <= a[126] * b[13] + a[127] * b[27] + a[128] * b[41] + a[129] * b[55] + a[130] * b[69] + a[131] * b[83] + a[132] * b[97] + a[133] * b[111] + a[134] * b[125] + a[135] * b[139] + a[136] * b[153] + a[137] * b[167] + a[138] * b[181] + a[139] * b[195];
                    c[140] <= a[140] * b[0] + a[141] * b[14] + a[142] * b[28] + a[143] * b[42] + a[144] * b[56] + a[145] * b[70] + a[146] * b[84] + a[147] * b[98] + a[148] * b[112] + a[149] * b[126] + a[150] * b[140] + a[151] * b[154] + a[152] * b[168] + a[153] * b[182];
                    c[141] <= a[140] * b[1] + a[141] * b[15] + a[142] * b[29] + a[143] * b[43] + a[144] * b[57] + a[145] * b[71] + a[146] * b[85] + a[147] * b[99] + a[148] * b[113] + a[149] * b[127] + a[150] * b[141] + a[151] * b[155] + a[152] * b[169] + a[153] * b[183];
                    c[142] <= a[140] * b[2] + a[141] * b[16] + a[142] * b[30] + a[143] * b[44] + a[144] * b[58] + a[145] * b[72] + a[146] * b[86] + a[147] * b[100] + a[148] * b[114] + a[149] * b[128] + a[150] * b[142] + a[151] * b[156] + a[152] * b[170] + a[153] * b[184];
                    c[143] <= a[140] * b[3] + a[141] * b[17] + a[142] * b[31] + a[143] * b[45] + a[144] * b[59] + a[145] * b[73] + a[146] * b[87] + a[147] * b[101] + a[148] * b[115] + a[149] * b[129] + a[150] * b[143] + a[151] * b[157] + a[152] * b[171] + a[153] * b[185];
                    c[144] <= a[140] * b[4] + a[141] * b[18] + a[142] * b[32] + a[143] * b[46] + a[144] * b[60] + a[145] * b[74] + a[146] * b[88] + a[147] * b[102] + a[148] * b[116] + a[149] * b[130] + a[150] * b[144] + a[151] * b[158] + a[152] * b[172] + a[153] * b[186];
                    c[145] <= a[140] * b[5] + a[141] * b[19] + a[142] * b[33] + a[143] * b[47] + a[144] * b[61] + a[145] * b[75] + a[146] * b[89] + a[147] * b[103] + a[148] * b[117] + a[149] * b[131] + a[150] * b[145] + a[151] * b[159] + a[152] * b[173] + a[153] * b[187];
                    c[146] <= a[140] * b[6] + a[141] * b[20] + a[142] * b[34] + a[143] * b[48] + a[144] * b[62] + a[145] * b[76] + a[146] * b[90] + a[147] * b[104] + a[148] * b[118] + a[149] * b[132] + a[150] * b[146] + a[151] * b[160] + a[152] * b[174] + a[153] * b[188];
                    c[147] <= a[140] * b[7] + a[141] * b[21] + a[142] * b[35] + a[143] * b[49] + a[144] * b[63] + a[145] * b[77] + a[146] * b[91] + a[147] * b[105] + a[148] * b[119] + a[149] * b[133] + a[150] * b[147] + a[151] * b[161] + a[152] * b[175] + a[153] * b[189];
                    c[148] <= a[140] * b[8] + a[141] * b[22] + a[142] * b[36] + a[143] * b[50] + a[144] * b[64] + a[145] * b[78] + a[146] * b[92] + a[147] * b[106] + a[148] * b[120] + a[149] * b[134] + a[150] * b[148] + a[151] * b[162] + a[152] * b[176] + a[153] * b[190];
                    c[149] <= a[140] * b[9] + a[141] * b[23] + a[142] * b[37] + a[143] * b[51] + a[144] * b[65] + a[145] * b[79] + a[146] * b[93] + a[147] * b[107] + a[148] * b[121] + a[149] * b[135] + a[150] * b[149] + a[151] * b[163] + a[152] * b[177] + a[153] * b[191];
                    c[150] <= a[140] * b[10] + a[141] * b[24] + a[142] * b[38] + a[143] * b[52] + a[144] * b[66] + a[145] * b[80] + a[146] * b[94] + a[147] * b[108] + a[148] * b[122] + a[149] * b[136] + a[150] * b[150] + a[151] * b[164] + a[152] * b[178] + a[153] * b[192];
                    c[151] <= a[140] * b[11] + a[141] * b[25] + a[142] * b[39] + a[143] * b[53] + a[144] * b[67] + a[145] * b[81] + a[146] * b[95] + a[147] * b[109] + a[148] * b[123] + a[149] * b[137] + a[150] * b[151] + a[151] * b[165] + a[152] * b[179] + a[153] * b[193];
                    c[152] <= a[140] * b[12] + a[141] * b[26] + a[142] * b[40] + a[143] * b[54] + a[144] * b[68] + a[145] * b[82] + a[146] * b[96] + a[147] * b[110] + a[148] * b[124] + a[149] * b[138] + a[150] * b[152] + a[151] * b[166] + a[152] * b[180] + a[153] * b[194];
                    c[153] <= a[140] * b[13] + a[141] * b[27] + a[142] * b[41] + a[143] * b[55] + a[144] * b[69] + a[145] * b[83] + a[146] * b[97] + a[147] * b[111] + a[148] * b[125] + a[149] * b[139] + a[150] * b[153] + a[151] * b[167] + a[152] * b[181] + a[153] * b[195];
                    c[154] <= a[154] * b[0] + a[155] * b[14] + a[156] * b[28] + a[157] * b[42] + a[158] * b[56] + a[159] * b[70] + a[160] * b[84] + a[161] * b[98] + a[162] * b[112] + a[163] * b[126] + a[164] * b[140] + a[165] * b[154] + a[166] * b[168] + a[167] * b[182];
                    c[155] <= a[154] * b[1] + a[155] * b[15] + a[156] * b[29] + a[157] * b[43] + a[158] * b[57] + a[159] * b[71] + a[160] * b[85] + a[161] * b[99] + a[162] * b[113] + a[163] * b[127] + a[164] * b[141] + a[165] * b[155] + a[166] * b[169] + a[167] * b[183];
                    c[156] <= a[154] * b[2] + a[155] * b[16] + a[156] * b[30] + a[157] * b[44] + a[158] * b[58] + a[159] * b[72] + a[160] * b[86] + a[161] * b[100] + a[162] * b[114] + a[163] * b[128] + a[164] * b[142] + a[165] * b[156] + a[166] * b[170] + a[167] * b[184];
                    c[157] <= a[154] * b[3] + a[155] * b[17] + a[156] * b[31] + a[157] * b[45] + a[158] * b[59] + a[159] * b[73] + a[160] * b[87] + a[161] * b[101] + a[162] * b[115] + a[163] * b[129] + a[164] * b[143] + a[165] * b[157] + a[166] * b[171] + a[167] * b[185];
                    c[158] <= a[154] * b[4] + a[155] * b[18] + a[156] * b[32] + a[157] * b[46] + a[158] * b[60] + a[159] * b[74] + a[160] * b[88] + a[161] * b[102] + a[162] * b[116] + a[163] * b[130] + a[164] * b[144] + a[165] * b[158] + a[166] * b[172] + a[167] * b[186];
                    c[159] <= a[154] * b[5] + a[155] * b[19] + a[156] * b[33] + a[157] * b[47] + a[158] * b[61] + a[159] * b[75] + a[160] * b[89] + a[161] * b[103] + a[162] * b[117] + a[163] * b[131] + a[164] * b[145] + a[165] * b[159] + a[166] * b[173] + a[167] * b[187];
                    c[160] <= a[154] * b[6] + a[155] * b[20] + a[156] * b[34] + a[157] * b[48] + a[158] * b[62] + a[159] * b[76] + a[160] * b[90] + a[161] * b[104] + a[162] * b[118] + a[163] * b[132] + a[164] * b[146] + a[165] * b[160] + a[166] * b[174] + a[167] * b[188];
                    c[161] <= a[154] * b[7] + a[155] * b[21] + a[156] * b[35] + a[157] * b[49] + a[158] * b[63] + a[159] * b[77] + a[160] * b[91] + a[161] * b[105] + a[162] * b[119] + a[163] * b[133] + a[164] * b[147] + a[165] * b[161] + a[166] * b[175] + a[167] * b[189];
                    c[162] <= a[154] * b[8] + a[155] * b[22] + a[156] * b[36] + a[157] * b[50] + a[158] * b[64] + a[159] * b[78] + a[160] * b[92] + a[161] * b[106] + a[162] * b[120] + a[163] * b[134] + a[164] * b[148] + a[165] * b[162] + a[166] * b[176] + a[167] * b[190];
                    c[163] <= a[154] * b[9] + a[155] * b[23] + a[156] * b[37] + a[157] * b[51] + a[158] * b[65] + a[159] * b[79] + a[160] * b[93] + a[161] * b[107] + a[162] * b[121] + a[163] * b[135] + a[164] * b[149] + a[165] * b[163] + a[166] * b[177] + a[167] * b[191];
                    c[164] <= a[154] * b[10] + a[155] * b[24] + a[156] * b[38] + a[157] * b[52] + a[158] * b[66] + a[159] * b[80] + a[160] * b[94] + a[161] * b[108] + a[162] * b[122] + a[163] * b[136] + a[164] * b[150] + a[165] * b[164] + a[166] * b[178] + a[167] * b[192];
                    c[165] <= a[154] * b[11] + a[155] * b[25] + a[156] * b[39] + a[157] * b[53] + a[158] * b[67] + a[159] * b[81] + a[160] * b[95] + a[161] * b[109] + a[162] * b[123] + a[163] * b[137] + a[164] * b[151] + a[165] * b[165] + a[166] * b[179] + a[167] * b[193];
                    c[166] <= a[154] * b[12] + a[155] * b[26] + a[156] * b[40] + a[157] * b[54] + a[158] * b[68] + a[159] * b[82] + a[160] * b[96] + a[161] * b[110] + a[162] * b[124] + a[163] * b[138] + a[164] * b[152] + a[165] * b[166] + a[166] * b[180] + a[167] * b[194];
                    c[167] <= a[154] * b[13] + a[155] * b[27] + a[156] * b[41] + a[157] * b[55] + a[158] * b[69] + a[159] * b[83] + a[160] * b[97] + a[161] * b[111] + a[162] * b[125] + a[163] * b[139] + a[164] * b[153] + a[165] * b[167] + a[166] * b[181] + a[167] * b[195];
                    c[168] <= a[168] * b[0] + a[169] * b[14] + a[170] * b[28] + a[171] * b[42] + a[172] * b[56] + a[173] * b[70] + a[174] * b[84] + a[175] * b[98] + a[176] * b[112] + a[177] * b[126] + a[178] * b[140] + a[179] * b[154] + a[180] * b[168] + a[181] * b[182];
                    c[169] <= a[168] * b[1] + a[169] * b[15] + a[170] * b[29] + a[171] * b[43] + a[172] * b[57] + a[173] * b[71] + a[174] * b[85] + a[175] * b[99] + a[176] * b[113] + a[177] * b[127] + a[178] * b[141] + a[179] * b[155] + a[180] * b[169] + a[181] * b[183];
                    c[170] <= a[168] * b[2] + a[169] * b[16] + a[170] * b[30] + a[171] * b[44] + a[172] * b[58] + a[173] * b[72] + a[174] * b[86] + a[175] * b[100] + a[176] * b[114] + a[177] * b[128] + a[178] * b[142] + a[179] * b[156] + a[180] * b[170] + a[181] * b[184];
                    c[171] <= a[168] * b[3] + a[169] * b[17] + a[170] * b[31] + a[171] * b[45] + a[172] * b[59] + a[173] * b[73] + a[174] * b[87] + a[175] * b[101] + a[176] * b[115] + a[177] * b[129] + a[178] * b[143] + a[179] * b[157] + a[180] * b[171] + a[181] * b[185];
                    c[172] <= a[168] * b[4] + a[169] * b[18] + a[170] * b[32] + a[171] * b[46] + a[172] * b[60] + a[173] * b[74] + a[174] * b[88] + a[175] * b[102] + a[176] * b[116] + a[177] * b[130] + a[178] * b[144] + a[179] * b[158] + a[180] * b[172] + a[181] * b[186];
                    c[173] <= a[168] * b[5] + a[169] * b[19] + a[170] * b[33] + a[171] * b[47] + a[172] * b[61] + a[173] * b[75] + a[174] * b[89] + a[175] * b[103] + a[176] * b[117] + a[177] * b[131] + a[178] * b[145] + a[179] * b[159] + a[180] * b[173] + a[181] * b[187];
                    c[174] <= a[168] * b[6] + a[169] * b[20] + a[170] * b[34] + a[171] * b[48] + a[172] * b[62] + a[173] * b[76] + a[174] * b[90] + a[175] * b[104] + a[176] * b[118] + a[177] * b[132] + a[178] * b[146] + a[179] * b[160] + a[180] * b[174] + a[181] * b[188];
                    c[175] <= a[168] * b[7] + a[169] * b[21] + a[170] * b[35] + a[171] * b[49] + a[172] * b[63] + a[173] * b[77] + a[174] * b[91] + a[175] * b[105] + a[176] * b[119] + a[177] * b[133] + a[178] * b[147] + a[179] * b[161] + a[180] * b[175] + a[181] * b[189];
                    c[176] <= a[168] * b[8] + a[169] * b[22] + a[170] * b[36] + a[171] * b[50] + a[172] * b[64] + a[173] * b[78] + a[174] * b[92] + a[175] * b[106] + a[176] * b[120] + a[177] * b[134] + a[178] * b[148] + a[179] * b[162] + a[180] * b[176] + a[181] * b[190];
                    c[177] <= a[168] * b[9] + a[169] * b[23] + a[170] * b[37] + a[171] * b[51] + a[172] * b[65] + a[173] * b[79] + a[174] * b[93] + a[175] * b[107] + a[176] * b[121] + a[177] * b[135] + a[178] * b[149] + a[179] * b[163] + a[180] * b[177] + a[181] * b[191];
                    c[178] <= a[168] * b[10] + a[169] * b[24] + a[170] * b[38] + a[171] * b[52] + a[172] * b[66] + a[173] * b[80] + a[174] * b[94] + a[175] * b[108] + a[176] * b[122] + a[177] * b[136] + a[178] * b[150] + a[179] * b[164] + a[180] * b[178] + a[181] * b[192];
                    c[179] <= a[168] * b[11] + a[169] * b[25] + a[170] * b[39] + a[171] * b[53] + a[172] * b[67] + a[173] * b[81] + a[174] * b[95] + a[175] * b[109] + a[176] * b[123] + a[177] * b[137] + a[178] * b[151] + a[179] * b[165] + a[180] * b[179] + a[181] * b[193];
                    c[180] <= a[168] * b[12] + a[169] * b[26] + a[170] * b[40] + a[171] * b[54] + a[172] * b[68] + a[173] * b[82] + a[174] * b[96] + a[175] * b[110] + a[176] * b[124] + a[177] * b[138] + a[178] * b[152] + a[179] * b[166] + a[180] * b[180] + a[181] * b[194];
                    c[181] <= a[168] * b[13] + a[169] * b[27] + a[170] * b[41] + a[171] * b[55] + a[172] * b[69] + a[173] * b[83] + a[174] * b[97] + a[175] * b[111] + a[176] * b[125] + a[177] * b[139] + a[178] * b[153] + a[179] * b[167] + a[180] * b[181] + a[181] * b[195];
                    c[182] <= a[182] * b[0] + a[183] * b[14] + a[184] * b[28] + a[185] * b[42] + a[186] * b[56] + a[187] * b[70] + a[188] * b[84] + a[189] * b[98] + a[190] * b[112] + a[191] * b[126] + a[192] * b[140] + a[193] * b[154] + a[194] * b[168] + a[195] * b[182];
                    c[183] <= a[182] * b[1] + a[183] * b[15] + a[184] * b[29] + a[185] * b[43] + a[186] * b[57] + a[187] * b[71] + a[188] * b[85] + a[189] * b[99] + a[190] * b[113] + a[191] * b[127] + a[192] * b[141] + a[193] * b[155] + a[194] * b[169] + a[195] * b[183];
                    c[184] <= a[182] * b[2] + a[183] * b[16] + a[184] * b[30] + a[185] * b[44] + a[186] * b[58] + a[187] * b[72] + a[188] * b[86] + a[189] * b[100] + a[190] * b[114] + a[191] * b[128] + a[192] * b[142] + a[193] * b[156] + a[194] * b[170] + a[195] * b[184];
                    c[185] <= a[182] * b[3] + a[183] * b[17] + a[184] * b[31] + a[185] * b[45] + a[186] * b[59] + a[187] * b[73] + a[188] * b[87] + a[189] * b[101] + a[190] * b[115] + a[191] * b[129] + a[192] * b[143] + a[193] * b[157] + a[194] * b[171] + a[195] * b[185];
                    c[186] <= a[182] * b[4] + a[183] * b[18] + a[184] * b[32] + a[185] * b[46] + a[186] * b[60] + a[187] * b[74] + a[188] * b[88] + a[189] * b[102] + a[190] * b[116] + a[191] * b[130] + a[192] * b[144] + a[193] * b[158] + a[194] * b[172] + a[195] * b[186];
                    c[187] <= a[182] * b[5] + a[183] * b[19] + a[184] * b[33] + a[185] * b[47] + a[186] * b[61] + a[187] * b[75] + a[188] * b[89] + a[189] * b[103] + a[190] * b[117] + a[191] * b[131] + a[192] * b[145] + a[193] * b[159] + a[194] * b[173] + a[195] * b[187];
                    c[188] <= a[182] * b[6] + a[183] * b[20] + a[184] * b[34] + a[185] * b[48] + a[186] * b[62] + a[187] * b[76] + a[188] * b[90] + a[189] * b[104] + a[190] * b[118] + a[191] * b[132] + a[192] * b[146] + a[193] * b[160] + a[194] * b[174] + a[195] * b[188];
                    c[189] <= a[182] * b[7] + a[183] * b[21] + a[184] * b[35] + a[185] * b[49] + a[186] * b[63] + a[187] * b[77] + a[188] * b[91] + a[189] * b[105] + a[190] * b[119] + a[191] * b[133] + a[192] * b[147] + a[193] * b[161] + a[194] * b[175] + a[195] * b[189];
                    c[190] <= a[182] * b[8] + a[183] * b[22] + a[184] * b[36] + a[185] * b[50] + a[186] * b[64] + a[187] * b[78] + a[188] * b[92] + a[189] * b[106] + a[190] * b[120] + a[191] * b[134] + a[192] * b[148] + a[193] * b[162] + a[194] * b[176] + a[195] * b[190];
                    c[191] <= a[182] * b[9] + a[183] * b[23] + a[184] * b[37] + a[185] * b[51] + a[186] * b[65] + a[187] * b[79] + a[188] * b[93] + a[189] * b[107] + a[190] * b[121] + a[191] * b[135] + a[192] * b[149] + a[193] * b[163] + a[194] * b[177] + a[195] * b[191];
                    c[192] <= a[182] * b[10] + a[183] * b[24] + a[184] * b[38] + a[185] * b[52] + a[186] * b[66] + a[187] * b[80] + a[188] * b[94] + a[189] * b[108] + a[190] * b[122] + a[191] * b[136] + a[192] * b[150] + a[193] * b[164] + a[194] * b[178] + a[195] * b[192];
                    c[193] <= a[182] * b[11] + a[183] * b[25] + a[184] * b[39] + a[185] * b[53] + a[186] * b[67] + a[187] * b[81] + a[188] * b[95] + a[189] * b[109] + a[190] * b[123] + a[191] * b[137] + a[192] * b[151] + a[193] * b[165] + a[194] * b[179] + a[195] * b[193];
                    c[194] <= a[182] * b[12] + a[183] * b[26] + a[184] * b[40] + a[185] * b[54] + a[186] * b[68] + a[187] * b[82] + a[188] * b[96] + a[189] * b[110] + a[190] * b[124] + a[191] * b[138] + a[192] * b[152] + a[193] * b[166] + a[194] * b[180] + a[195] * b[194];
                    c[195] <= a[182] * b[13] + a[183] * b[27] + a[184] * b[41] + a[185] * b[55] + a[186] * b[69] + a[187] * b[83] + a[188] * b[97] + a[189] * b[111] + a[190] * b[125] + a[191] * b[139] + a[192] * b[153] + a[193] * b[167] + a[194] * b[181] + a[195] * b[195];
                    c[196] <= a[196] * b[0] + a[197] * b[14] + a[198] * b[28] + a[199] * b[42] + a[200] * b[56] + a[201] * b[70] + a[202] * b[84] + a[203] * b[98] + a[204] * b[112] + a[205] * b[126] + a[206] * b[140] + a[207] * b[154] + a[208] * b[168] + a[209] * b[182];
                    c[197] <= a[196] * b[1] + a[197] * b[15] + a[198] * b[29] + a[199] * b[43] + a[200] * b[57] + a[201] * b[71] + a[202] * b[85] + a[203] * b[99] + a[204] * b[113] + a[205] * b[127] + a[206] * b[141] + a[207] * b[155] + a[208] * b[169] + a[209] * b[183];
                    c[198] <= a[196] * b[2] + a[197] * b[16] + a[198] * b[30] + a[199] * b[44] + a[200] * b[58] + a[201] * b[72] + a[202] * b[86] + a[203] * b[100] + a[204] * b[114] + a[205] * b[128] + a[206] * b[142] + a[207] * b[156] + a[208] * b[170] + a[209] * b[184];
                    c[199] <= a[196] * b[3] + a[197] * b[17] + a[198] * b[31] + a[199] * b[45] + a[200] * b[59] + a[201] * b[73] + a[202] * b[87] + a[203] * b[101] + a[204] * b[115] + a[205] * b[129] + a[206] * b[143] + a[207] * b[157] + a[208] * b[171] + a[209] * b[185];
                    c[200] <= a[196] * b[4] + a[197] * b[18] + a[198] * b[32] + a[199] * b[46] + a[200] * b[60] + a[201] * b[74] + a[202] * b[88] + a[203] * b[102] + a[204] * b[116] + a[205] * b[130] + a[206] * b[144] + a[207] * b[158] + a[208] * b[172] + a[209] * b[186];
                    c[201] <= a[196] * b[5] + a[197] * b[19] + a[198] * b[33] + a[199] * b[47] + a[200] * b[61] + a[201] * b[75] + a[202] * b[89] + a[203] * b[103] + a[204] * b[117] + a[205] * b[131] + a[206] * b[145] + a[207] * b[159] + a[208] * b[173] + a[209] * b[187];
                    c[202] <= a[196] * b[6] + a[197] * b[20] + a[198] * b[34] + a[199] * b[48] + a[200] * b[62] + a[201] * b[76] + a[202] * b[90] + a[203] * b[104] + a[204] * b[118] + a[205] * b[132] + a[206] * b[146] + a[207] * b[160] + a[208] * b[174] + a[209] * b[188];
                    c[203] <= a[196] * b[7] + a[197] * b[21] + a[198] * b[35] + a[199] * b[49] + a[200] * b[63] + a[201] * b[77] + a[202] * b[91] + a[203] * b[105] + a[204] * b[119] + a[205] * b[133] + a[206] * b[147] + a[207] * b[161] + a[208] * b[175] + a[209] * b[189];
                    c[204] <= a[196] * b[8] + a[197] * b[22] + a[198] * b[36] + a[199] * b[50] + a[200] * b[64] + a[201] * b[78] + a[202] * b[92] + a[203] * b[106] + a[204] * b[120] + a[205] * b[134] + a[206] * b[148] + a[207] * b[162] + a[208] * b[176] + a[209] * b[190];
                    c[205] <= a[196] * b[9] + a[197] * b[23] + a[198] * b[37] + a[199] * b[51] + a[200] * b[65] + a[201] * b[79] + a[202] * b[93] + a[203] * b[107] + a[204] * b[121] + a[205] * b[135] + a[206] * b[149] + a[207] * b[163] + a[208] * b[177] + a[209] * b[191];
                    c[206] <= a[196] * b[10] + a[197] * b[24] + a[198] * b[38] + a[199] * b[52] + a[200] * b[66] + a[201] * b[80] + a[202] * b[94] + a[203] * b[108] + a[204] * b[122] + a[205] * b[136] + a[206] * b[150] + a[207] * b[164] + a[208] * b[178] + a[209] * b[192];
                    c[207] <= a[196] * b[11] + a[197] * b[25] + a[198] * b[39] + a[199] * b[53] + a[200] * b[67] + a[201] * b[81] + a[202] * b[95] + a[203] * b[109] + a[204] * b[123] + a[205] * b[137] + a[206] * b[151] + a[207] * b[165] + a[208] * b[179] + a[209] * b[193];
                    c[208] <= a[196] * b[12] + a[197] * b[26] + a[198] * b[40] + a[199] * b[54] + a[200] * b[68] + a[201] * b[82] + a[202] * b[96] + a[203] * b[110] + a[204] * b[124] + a[205] * b[138] + a[206] * b[152] + a[207] * b[166] + a[208] * b[180] + a[209] * b[194];
                    c[209] <= a[196] * b[13] + a[197] * b[27] + a[198] * b[41] + a[199] * b[55] + a[200] * b[69] + a[201] * b[83] + a[202] * b[97] + a[203] * b[111] + a[204] * b[125] + a[205] * b[139] + a[206] * b[153] + a[207] * b[167] + a[208] * b[181] + a[209] * b[195];
                    c[210] <= a[210] * b[0] + a[211] * b[14] + a[212] * b[28] + a[213] * b[42] + a[214] * b[56] + a[215] * b[70] + a[216] * b[84] + a[217] * b[98] + a[218] * b[112] + a[219] * b[126] + a[220] * b[140] + a[221] * b[154] + a[222] * b[168] + a[223] * b[182];
                    c[211] <= a[210] * b[1] + a[211] * b[15] + a[212] * b[29] + a[213] * b[43] + a[214] * b[57] + a[215] * b[71] + a[216] * b[85] + a[217] * b[99] + a[218] * b[113] + a[219] * b[127] + a[220] * b[141] + a[221] * b[155] + a[222] * b[169] + a[223] * b[183];
                    c[212] <= a[210] * b[2] + a[211] * b[16] + a[212] * b[30] + a[213] * b[44] + a[214] * b[58] + a[215] * b[72] + a[216] * b[86] + a[217] * b[100] + a[218] * b[114] + a[219] * b[128] + a[220] * b[142] + a[221] * b[156] + a[222] * b[170] + a[223] * b[184];
                    c[213] <= a[210] * b[3] + a[211] * b[17] + a[212] * b[31] + a[213] * b[45] + a[214] * b[59] + a[215] * b[73] + a[216] * b[87] + a[217] * b[101] + a[218] * b[115] + a[219] * b[129] + a[220] * b[143] + a[221] * b[157] + a[222] * b[171] + a[223] * b[185];
                    c[214] <= a[210] * b[4] + a[211] * b[18] + a[212] * b[32] + a[213] * b[46] + a[214] * b[60] + a[215] * b[74] + a[216] * b[88] + a[217] * b[102] + a[218] * b[116] + a[219] * b[130] + a[220] * b[144] + a[221] * b[158] + a[222] * b[172] + a[223] * b[186];
                    c[215] <= a[210] * b[5] + a[211] * b[19] + a[212] * b[33] + a[213] * b[47] + a[214] * b[61] + a[215] * b[75] + a[216] * b[89] + a[217] * b[103] + a[218] * b[117] + a[219] * b[131] + a[220] * b[145] + a[221] * b[159] + a[222] * b[173] + a[223] * b[187];
                    c[216] <= a[210] * b[6] + a[211] * b[20] + a[212] * b[34] + a[213] * b[48] + a[214] * b[62] + a[215] * b[76] + a[216] * b[90] + a[217] * b[104] + a[218] * b[118] + a[219] * b[132] + a[220] * b[146] + a[221] * b[160] + a[222] * b[174] + a[223] * b[188];
                    c[217] <= a[210] * b[7] + a[211] * b[21] + a[212] * b[35] + a[213] * b[49] + a[214] * b[63] + a[215] * b[77] + a[216] * b[91] + a[217] * b[105] + a[218] * b[119] + a[219] * b[133] + a[220] * b[147] + a[221] * b[161] + a[222] * b[175] + a[223] * b[189];
                    c[218] <= a[210] * b[8] + a[211] * b[22] + a[212] * b[36] + a[213] * b[50] + a[214] * b[64] + a[215] * b[78] + a[216] * b[92] + a[217] * b[106] + a[218] * b[120] + a[219] * b[134] + a[220] * b[148] + a[221] * b[162] + a[222] * b[176] + a[223] * b[190];
                    c[219] <= a[210] * b[9] + a[211] * b[23] + a[212] * b[37] + a[213] * b[51] + a[214] * b[65] + a[215] * b[79] + a[216] * b[93] + a[217] * b[107] + a[218] * b[121] + a[219] * b[135] + a[220] * b[149] + a[221] * b[163] + a[222] * b[177] + a[223] * b[191];
                    c[220] <= a[210] * b[10] + a[211] * b[24] + a[212] * b[38] + a[213] * b[52] + a[214] * b[66] + a[215] * b[80] + a[216] * b[94] + a[217] * b[108] + a[218] * b[122] + a[219] * b[136] + a[220] * b[150] + a[221] * b[164] + a[222] * b[178] + a[223] * b[192];
                    c[221] <= a[210] * b[11] + a[211] * b[25] + a[212] * b[39] + a[213] * b[53] + a[214] * b[67] + a[215] * b[81] + a[216] * b[95] + a[217] * b[109] + a[218] * b[123] + a[219] * b[137] + a[220] * b[151] + a[221] * b[165] + a[222] * b[179] + a[223] * b[193];
                    c[222] <= a[210] * b[12] + a[211] * b[26] + a[212] * b[40] + a[213] * b[54] + a[214] * b[68] + a[215] * b[82] + a[216] * b[96] + a[217] * b[110] + a[218] * b[124] + a[219] * b[138] + a[220] * b[152] + a[221] * b[166] + a[222] * b[180] + a[223] * b[194];
                    c[223] <= a[210] * b[13] + a[211] * b[27] + a[212] * b[41] + a[213] * b[55] + a[214] * b[69] + a[215] * b[83] + a[216] * b[97] + a[217] * b[111] + a[218] * b[125] + a[219] * b[139] + a[220] * b[153] + a[221] * b[167] + a[222] * b[181] + a[223] * b[195];
                    c[224] <= a[224] * b[0] + a[225] * b[14] + a[226] * b[28] + a[227] * b[42] + a[228] * b[56] + a[229] * b[70] + a[230] * b[84] + a[231] * b[98] + a[232] * b[112] + a[233] * b[126] + a[234] * b[140] + a[235] * b[154] + a[236] * b[168] + a[237] * b[182];
                    c[225] <= a[224] * b[1] + a[225] * b[15] + a[226] * b[29] + a[227] * b[43] + a[228] * b[57] + a[229] * b[71] + a[230] * b[85] + a[231] * b[99] + a[232] * b[113] + a[233] * b[127] + a[234] * b[141] + a[235] * b[155] + a[236] * b[169] + a[237] * b[183];
                    c[226] <= a[224] * b[2] + a[225] * b[16] + a[226] * b[30] + a[227] * b[44] + a[228] * b[58] + a[229] * b[72] + a[230] * b[86] + a[231] * b[100] + a[232] * b[114] + a[233] * b[128] + a[234] * b[142] + a[235] * b[156] + a[236] * b[170] + a[237] * b[184];
                    c[227] <= a[224] * b[3] + a[225] * b[17] + a[226] * b[31] + a[227] * b[45] + a[228] * b[59] + a[229] * b[73] + a[230] * b[87] + a[231] * b[101] + a[232] * b[115] + a[233] * b[129] + a[234] * b[143] + a[235] * b[157] + a[236] * b[171] + a[237] * b[185];
                    c[228] <= a[224] * b[4] + a[225] * b[18] + a[226] * b[32] + a[227] * b[46] + a[228] * b[60] + a[229] * b[74] + a[230] * b[88] + a[231] * b[102] + a[232] * b[116] + a[233] * b[130] + a[234] * b[144] + a[235] * b[158] + a[236] * b[172] + a[237] * b[186];
                    c[229] <= a[224] * b[5] + a[225] * b[19] + a[226] * b[33] + a[227] * b[47] + a[228] * b[61] + a[229] * b[75] + a[230] * b[89] + a[231] * b[103] + a[232] * b[117] + a[233] * b[131] + a[234] * b[145] + a[235] * b[159] + a[236] * b[173] + a[237] * b[187];
                    c[230] <= a[224] * b[6] + a[225] * b[20] + a[226] * b[34] + a[227] * b[48] + a[228] * b[62] + a[229] * b[76] + a[230] * b[90] + a[231] * b[104] + a[232] * b[118] + a[233] * b[132] + a[234] * b[146] + a[235] * b[160] + a[236] * b[174] + a[237] * b[188];
                    c[231] <= a[224] * b[7] + a[225] * b[21] + a[226] * b[35] + a[227] * b[49] + a[228] * b[63] + a[229] * b[77] + a[230] * b[91] + a[231] * b[105] + a[232] * b[119] + a[233] * b[133] + a[234] * b[147] + a[235] * b[161] + a[236] * b[175] + a[237] * b[189];
                    c[232] <= a[224] * b[8] + a[225] * b[22] + a[226] * b[36] + a[227] * b[50] + a[228] * b[64] + a[229] * b[78] + a[230] * b[92] + a[231] * b[106] + a[232] * b[120] + a[233] * b[134] + a[234] * b[148] + a[235] * b[162] + a[236] * b[176] + a[237] * b[190];
                    c[233] <= a[224] * b[9] + a[225] * b[23] + a[226] * b[37] + a[227] * b[51] + a[228] * b[65] + a[229] * b[79] + a[230] * b[93] + a[231] * b[107] + a[232] * b[121] + a[233] * b[135] + a[234] * b[149] + a[235] * b[163] + a[236] * b[177] + a[237] * b[191];
                    c[234] <= a[224] * b[10] + a[225] * b[24] + a[226] * b[38] + a[227] * b[52] + a[228] * b[66] + a[229] * b[80] + a[230] * b[94] + a[231] * b[108] + a[232] * b[122] + a[233] * b[136] + a[234] * b[150] + a[235] * b[164] + a[236] * b[178] + a[237] * b[192];
                    c[235] <= a[224] * b[11] + a[225] * b[25] + a[226] * b[39] + a[227] * b[53] + a[228] * b[67] + a[229] * b[81] + a[230] * b[95] + a[231] * b[109] + a[232] * b[123] + a[233] * b[137] + a[234] * b[151] + a[235] * b[165] + a[236] * b[179] + a[237] * b[193];
                    c[236] <= a[224] * b[12] + a[225] * b[26] + a[226] * b[40] + a[227] * b[54] + a[228] * b[68] + a[229] * b[82] + a[230] * b[96] + a[231] * b[110] + a[232] * b[124] + a[233] * b[138] + a[234] * b[152] + a[235] * b[166] + a[236] * b[180] + a[237] * b[194];
                    c[237] <= a[224] * b[13] + a[225] * b[27] + a[226] * b[41] + a[227] * b[55] + a[228] * b[69] + a[229] * b[83] + a[230] * b[97] + a[231] * b[111] + a[232] * b[125] + a[233] * b[139] + a[234] * b[153] + a[235] * b[167] + a[236] * b[181] + a[237] * b[195];
                    c[238] <= a[238] * b[0] + a[239] * b[14] + a[240] * b[28] + a[241] * b[42] + a[242] * b[56] + a[243] * b[70] + a[244] * b[84] + a[245] * b[98] + a[246] * b[112] + a[247] * b[126] + a[248] * b[140] + a[249] * b[154] + a[250] * b[168] + a[251] * b[182];
                    c[239] <= a[238] * b[1] + a[239] * b[15] + a[240] * b[29] + a[241] * b[43] + a[242] * b[57] + a[243] * b[71] + a[244] * b[85] + a[245] * b[99] + a[246] * b[113] + a[247] * b[127] + a[248] * b[141] + a[249] * b[155] + a[250] * b[169] + a[251] * b[183];
                    c[240] <= a[238] * b[2] + a[239] * b[16] + a[240] * b[30] + a[241] * b[44] + a[242] * b[58] + a[243] * b[72] + a[244] * b[86] + a[245] * b[100] + a[246] * b[114] + a[247] * b[128] + a[248] * b[142] + a[249] * b[156] + a[250] * b[170] + a[251] * b[184];
                    c[241] <= a[238] * b[3] + a[239] * b[17] + a[240] * b[31] + a[241] * b[45] + a[242] * b[59] + a[243] * b[73] + a[244] * b[87] + a[245] * b[101] + a[246] * b[115] + a[247] * b[129] + a[248] * b[143] + a[249] * b[157] + a[250] * b[171] + a[251] * b[185];
                    c[242] <= a[238] * b[4] + a[239] * b[18] + a[240] * b[32] + a[241] * b[46] + a[242] * b[60] + a[243] * b[74] + a[244] * b[88] + a[245] * b[102] + a[246] * b[116] + a[247] * b[130] + a[248] * b[144] + a[249] * b[158] + a[250] * b[172] + a[251] * b[186];
                    c[243] <= a[238] * b[5] + a[239] * b[19] + a[240] * b[33] + a[241] * b[47] + a[242] * b[61] + a[243] * b[75] + a[244] * b[89] + a[245] * b[103] + a[246] * b[117] + a[247] * b[131] + a[248] * b[145] + a[249] * b[159] + a[250] * b[173] + a[251] * b[187];
                    c[244] <= a[238] * b[6] + a[239] * b[20] + a[240] * b[34] + a[241] * b[48] + a[242] * b[62] + a[243] * b[76] + a[244] * b[90] + a[245] * b[104] + a[246] * b[118] + a[247] * b[132] + a[248] * b[146] + a[249] * b[160] + a[250] * b[174] + a[251] * b[188];
                    c[245] <= a[238] * b[7] + a[239] * b[21] + a[240] * b[35] + a[241] * b[49] + a[242] * b[63] + a[243] * b[77] + a[244] * b[91] + a[245] * b[105] + a[246] * b[119] + a[247] * b[133] + a[248] * b[147] + a[249] * b[161] + a[250] * b[175] + a[251] * b[189];
                    c[246] <= a[238] * b[8] + a[239] * b[22] + a[240] * b[36] + a[241] * b[50] + a[242] * b[64] + a[243] * b[78] + a[244] * b[92] + a[245] * b[106] + a[246] * b[120] + a[247] * b[134] + a[248] * b[148] + a[249] * b[162] + a[250] * b[176] + a[251] * b[190];
                    c[247] <= a[238] * b[9] + a[239] * b[23] + a[240] * b[37] + a[241] * b[51] + a[242] * b[65] + a[243] * b[79] + a[244] * b[93] + a[245] * b[107] + a[246] * b[121] + a[247] * b[135] + a[248] * b[149] + a[249] * b[163] + a[250] * b[177] + a[251] * b[191];
                    c[248] <= a[238] * b[10] + a[239] * b[24] + a[240] * b[38] + a[241] * b[52] + a[242] * b[66] + a[243] * b[80] + a[244] * b[94] + a[245] * b[108] + a[246] * b[122] + a[247] * b[136] + a[248] * b[150] + a[249] * b[164] + a[250] * b[178] + a[251] * b[192];
                    c[249] <= a[238] * b[11] + a[239] * b[25] + a[240] * b[39] + a[241] * b[53] + a[242] * b[67] + a[243] * b[81] + a[244] * b[95] + a[245] * b[109] + a[246] * b[123] + a[247] * b[137] + a[248] * b[151] + a[249] * b[165] + a[250] * b[179] + a[251] * b[193];
                    c[250] <= a[238] * b[12] + a[239] * b[26] + a[240] * b[40] + a[241] * b[54] + a[242] * b[68] + a[243] * b[82] + a[244] * b[96] + a[245] * b[110] + a[246] * b[124] + a[247] * b[138] + a[248] * b[152] + a[249] * b[166] + a[250] * b[180] + a[251] * b[194];
                    c[251] <= a[238] * b[13] + a[239] * b[27] + a[240] * b[41] + a[241] * b[55] + a[242] * b[69] + a[243] * b[83] + a[244] * b[97] + a[245] * b[111] + a[246] * b[125] + a[247] * b[139] + a[248] * b[153] + a[249] * b[167] + a[250] * b[181] + a[251] * b[195];
                    c[252] <= a[252] * b[0] + a[253] * b[14] + a[254] * b[28] + a[255] * b[42] + a[256] * b[56] + a[257] * b[70] + a[258] * b[84] + a[259] * b[98] + a[260] * b[112] + a[261] * b[126] + a[262] * b[140] + a[263] * b[154] + a[264] * b[168] + a[265] * b[182];
                    c[253] <= a[252] * b[1] + a[253] * b[15] + a[254] * b[29] + a[255] * b[43] + a[256] * b[57] + a[257] * b[71] + a[258] * b[85] + a[259] * b[99] + a[260] * b[113] + a[261] * b[127] + a[262] * b[141] + a[263] * b[155] + a[264] * b[169] + a[265] * b[183];
                    c[254] <= a[252] * b[2] + a[253] * b[16] + a[254] * b[30] + a[255] * b[44] + a[256] * b[58] + a[257] * b[72] + a[258] * b[86] + a[259] * b[100] + a[260] * b[114] + a[261] * b[128] + a[262] * b[142] + a[263] * b[156] + a[264] * b[170] + a[265] * b[184];
                    c[255] <= a[252] * b[3] + a[253] * b[17] + a[254] * b[31] + a[255] * b[45] + a[256] * b[59] + a[257] * b[73] + a[258] * b[87] + a[259] * b[101] + a[260] * b[115] + a[261] * b[129] + a[262] * b[143] + a[263] * b[157] + a[264] * b[171] + a[265] * b[185];
                    c[256] <= a[252] * b[4] + a[253] * b[18] + a[254] * b[32] + a[255] * b[46] + a[256] * b[60] + a[257] * b[74] + a[258] * b[88] + a[259] * b[102] + a[260] * b[116] + a[261] * b[130] + a[262] * b[144] + a[263] * b[158] + a[264] * b[172] + a[265] * b[186];
                    c[257] <= a[252] * b[5] + a[253] * b[19] + a[254] * b[33] + a[255] * b[47] + a[256] * b[61] + a[257] * b[75] + a[258] * b[89] + a[259] * b[103] + a[260] * b[117] + a[261] * b[131] + a[262] * b[145] + a[263] * b[159] + a[264] * b[173] + a[265] * b[187];
                    c[258] <= a[252] * b[6] + a[253] * b[20] + a[254] * b[34] + a[255] * b[48] + a[256] * b[62] + a[257] * b[76] + a[258] * b[90] + a[259] * b[104] + a[260] * b[118] + a[261] * b[132] + a[262] * b[146] + a[263] * b[160] + a[264] * b[174] + a[265] * b[188];
                    c[259] <= a[252] * b[7] + a[253] * b[21] + a[254] * b[35] + a[255] * b[49] + a[256] * b[63] + a[257] * b[77] + a[258] * b[91] + a[259] * b[105] + a[260] * b[119] + a[261] * b[133] + a[262] * b[147] + a[263] * b[161] + a[264] * b[175] + a[265] * b[189];
                    c[260] <= a[252] * b[8] + a[253] * b[22] + a[254] * b[36] + a[255] * b[50] + a[256] * b[64] + a[257] * b[78] + a[258] * b[92] + a[259] * b[106] + a[260] * b[120] + a[261] * b[134] + a[262] * b[148] + a[263] * b[162] + a[264] * b[176] + a[265] * b[190];
                    c[261] <= a[252] * b[9] + a[253] * b[23] + a[254] * b[37] + a[255] * b[51] + a[256] * b[65] + a[257] * b[79] + a[258] * b[93] + a[259] * b[107] + a[260] * b[121] + a[261] * b[135] + a[262] * b[149] + a[263] * b[163] + a[264] * b[177] + a[265] * b[191];
                    c[262] <= a[252] * b[10] + a[253] * b[24] + a[254] * b[38] + a[255] * b[52] + a[256] * b[66] + a[257] * b[80] + a[258] * b[94] + a[259] * b[108] + a[260] * b[122] + a[261] * b[136] + a[262] * b[150] + a[263] * b[164] + a[264] * b[178] + a[265] * b[192];
                    c[263] <= a[252] * b[11] + a[253] * b[25] + a[254] * b[39] + a[255] * b[53] + a[256] * b[67] + a[257] * b[81] + a[258] * b[95] + a[259] * b[109] + a[260] * b[123] + a[261] * b[137] + a[262] * b[151] + a[263] * b[165] + a[264] * b[179] + a[265] * b[193];
                    c[264] <= a[252] * b[12] + a[253] * b[26] + a[254] * b[40] + a[255] * b[54] + a[256] * b[68] + a[257] * b[82] + a[258] * b[96] + a[259] * b[110] + a[260] * b[124] + a[261] * b[138] + a[262] * b[152] + a[263] * b[166] + a[264] * b[180] + a[265] * b[194];
                    c[265] <= a[252] * b[13] + a[253] * b[27] + a[254] * b[41] + a[255] * b[55] + a[256] * b[69] + a[257] * b[83] + a[258] * b[97] + a[259] * b[111] + a[260] * b[125] + a[261] * b[139] + a[262] * b[153] + a[263] * b[167] + a[264] * b[181] + a[265] * b[195];
                    c[266] <= a[266] * b[0] + a[267] * b[14] + a[268] * b[28] + a[269] * b[42] + a[270] * b[56] + a[271] * b[70] + a[272] * b[84] + a[273] * b[98] + a[274] * b[112] + a[275] * b[126] + a[276] * b[140] + a[277] * b[154] + a[278] * b[168] + a[279] * b[182];
                    c[267] <= a[266] * b[1] + a[267] * b[15] + a[268] * b[29] + a[269] * b[43] + a[270] * b[57] + a[271] * b[71] + a[272] * b[85] + a[273] * b[99] + a[274] * b[113] + a[275] * b[127] + a[276] * b[141] + a[277] * b[155] + a[278] * b[169] + a[279] * b[183];
                    c[268] <= a[266] * b[2] + a[267] * b[16] + a[268] * b[30] + a[269] * b[44] + a[270] * b[58] + a[271] * b[72] + a[272] * b[86] + a[273] * b[100] + a[274] * b[114] + a[275] * b[128] + a[276] * b[142] + a[277] * b[156] + a[278] * b[170] + a[279] * b[184];
                    c[269] <= a[266] * b[3] + a[267] * b[17] + a[268] * b[31] + a[269] * b[45] + a[270] * b[59] + a[271] * b[73] + a[272] * b[87] + a[273] * b[101] + a[274] * b[115] + a[275] * b[129] + a[276] * b[143] + a[277] * b[157] + a[278] * b[171] + a[279] * b[185];
                    c[270] <= a[266] * b[4] + a[267] * b[18] + a[268] * b[32] + a[269] * b[46] + a[270] * b[60] + a[271] * b[74] + a[272] * b[88] + a[273] * b[102] + a[274] * b[116] + a[275] * b[130] + a[276] * b[144] + a[277] * b[158] + a[278] * b[172] + a[279] * b[186];
                    c[271] <= a[266] * b[5] + a[267] * b[19] + a[268] * b[33] + a[269] * b[47] + a[270] * b[61] + a[271] * b[75] + a[272] * b[89] + a[273] * b[103] + a[274] * b[117] + a[275] * b[131] + a[276] * b[145] + a[277] * b[159] + a[278] * b[173] + a[279] * b[187];
                    c[272] <= a[266] * b[6] + a[267] * b[20] + a[268] * b[34] + a[269] * b[48] + a[270] * b[62] + a[271] * b[76] + a[272] * b[90] + a[273] * b[104] + a[274] * b[118] + a[275] * b[132] + a[276] * b[146] + a[277] * b[160] + a[278] * b[174] + a[279] * b[188];
                    c[273] <= a[266] * b[7] + a[267] * b[21] + a[268] * b[35] + a[269] * b[49] + a[270] * b[63] + a[271] * b[77] + a[272] * b[91] + a[273] * b[105] + a[274] * b[119] + a[275] * b[133] + a[276] * b[147] + a[277] * b[161] + a[278] * b[175] + a[279] * b[189];
                    c[274] <= a[266] * b[8] + a[267] * b[22] + a[268] * b[36] + a[269] * b[50] + a[270] * b[64] + a[271] * b[78] + a[272] * b[92] + a[273] * b[106] + a[274] * b[120] + a[275] * b[134] + a[276] * b[148] + a[277] * b[162] + a[278] * b[176] + a[279] * b[190];
                    c[275] <= a[266] * b[9] + a[267] * b[23] + a[268] * b[37] + a[269] * b[51] + a[270] * b[65] + a[271] * b[79] + a[272] * b[93] + a[273] * b[107] + a[274] * b[121] + a[275] * b[135] + a[276] * b[149] + a[277] * b[163] + a[278] * b[177] + a[279] * b[191];
                    c[276] <= a[266] * b[10] + a[267] * b[24] + a[268] * b[38] + a[269] * b[52] + a[270] * b[66] + a[271] * b[80] + a[272] * b[94] + a[273] * b[108] + a[274] * b[122] + a[275] * b[136] + a[276] * b[150] + a[277] * b[164] + a[278] * b[178] + a[279] * b[192];
                    c[277] <= a[266] * b[11] + a[267] * b[25] + a[268] * b[39] + a[269] * b[53] + a[270] * b[67] + a[271] * b[81] + a[272] * b[95] + a[273] * b[109] + a[274] * b[123] + a[275] * b[137] + a[276] * b[151] + a[277] * b[165] + a[278] * b[179] + a[279] * b[193];
                    c[278] <= a[266] * b[12] + a[267] * b[26] + a[268] * b[40] + a[269] * b[54] + a[270] * b[68] + a[271] * b[82] + a[272] * b[96] + a[273] * b[110] + a[274] * b[124] + a[275] * b[138] + a[276] * b[152] + a[277] * b[166] + a[278] * b[180] + a[279] * b[194];
                    c[279] <= a[266] * b[13] + a[267] * b[27] + a[268] * b[41] + a[269] * b[55] + a[270] * b[69] + a[271] * b[83] + a[272] * b[97] + a[273] * b[111] + a[274] * b[125] + a[275] * b[139] + a[276] * b[153] + a[277] * b[167] + a[278] * b[181] + a[279] * b[195];
                end
            endcase
        end
    end

    always @(posedge clk) begin
        if (rst) begin
            state <= 0;
        end else begin
            case (state)
                fin: begin
                    if (matmult_accept) begin
                        state <= idle;
                    end
                end
                idle: begin
                    if (matmult_ready) begin
                        state <= calc;
                    end
                end
                calc: begin
                    state <= fin;
                end
            endcase
        end
    end

endmodule
