module listc20r14_matmult (
    input wire clk,
    input wire rst,
    input wire matmult_ready,
    input wire matmult_accept,
    output reg matmult_valid,
    input wire signed [63:0] matmult_in_a0,
    input wire signed [63:0] matmult_in_a1,
    input wire signed [63:0] matmult_in_a2,
    input wire signed [63:0] matmult_in_a3,
    input wire signed [63:0] matmult_in_a4,
    input wire signed [63:0] matmult_in_a5,
    input wire signed [63:0] matmult_in_a6,
    input wire signed [63:0] matmult_in_a7,
    input wire signed [63:0] matmult_in_a8,
    input wire signed [63:0] matmult_in_a9,
    input wire signed [63:0] matmult_in_a10,
    input wire signed [63:0] matmult_in_a11,
    input wire signed [63:0] matmult_in_a12,
    input wire signed [63:0] matmult_in_a13,
    input wire signed [63:0] matmult_in_a14,
    input wire signed [63:0] matmult_in_a15,
    input wire signed [63:0] matmult_in_a16,
    input wire signed [63:0] matmult_in_a17,
    input wire signed [63:0] matmult_in_a18,
    input wire signed [63:0] matmult_in_a19,
    input wire signed [63:0] matmult_in_a20,
    input wire signed [63:0] matmult_in_a21,
    input wire signed [63:0] matmult_in_a22,
    input wire signed [63:0] matmult_in_a23,
    input wire signed [63:0] matmult_in_a24,
    input wire signed [63:0] matmult_in_a25,
    input wire signed [63:0] matmult_in_a26,
    input wire signed [63:0] matmult_in_a27,
    input wire signed [63:0] matmult_in_a28,
    input wire signed [63:0] matmult_in_a29,
    input wire signed [63:0] matmult_in_a30,
    input wire signed [63:0] matmult_in_a31,
    input wire signed [63:0] matmult_in_a32,
    input wire signed [63:0] matmult_in_a33,
    input wire signed [63:0] matmult_in_a34,
    input wire signed [63:0] matmult_in_a35,
    input wire signed [63:0] matmult_in_a36,
    input wire signed [63:0] matmult_in_a37,
    input wire signed [63:0] matmult_in_a38,
    input wire signed [63:0] matmult_in_a39,
    input wire signed [63:0] matmult_in_a40,
    input wire signed [63:0] matmult_in_a41,
    input wire signed [63:0] matmult_in_a42,
    input wire signed [63:0] matmult_in_a43,
    input wire signed [63:0] matmult_in_a44,
    input wire signed [63:0] matmult_in_a45,
    input wire signed [63:0] matmult_in_a46,
    input wire signed [63:0] matmult_in_a47,
    input wire signed [63:0] matmult_in_a48,
    input wire signed [63:0] matmult_in_a49,
    input wire signed [63:0] matmult_in_a50,
    input wire signed [63:0] matmult_in_a51,
    input wire signed [63:0] matmult_in_a52,
    input wire signed [63:0] matmult_in_a53,
    input wire signed [63:0] matmult_in_a54,
    input wire signed [63:0] matmult_in_a55,
    input wire signed [63:0] matmult_in_a56,
    input wire signed [63:0] matmult_in_a57,
    input wire signed [63:0] matmult_in_a58,
    input wire signed [63:0] matmult_in_a59,
    input wire signed [63:0] matmult_in_a60,
    input wire signed [63:0] matmult_in_a61,
    input wire signed [63:0] matmult_in_a62,
    input wire signed [63:0] matmult_in_a63,
    input wire signed [63:0] matmult_in_a64,
    input wire signed [63:0] matmult_in_a65,
    input wire signed [63:0] matmult_in_a66,
    input wire signed [63:0] matmult_in_a67,
    input wire signed [63:0] matmult_in_a68,
    input wire signed [63:0] matmult_in_a69,
    input wire signed [63:0] matmult_in_a70,
    input wire signed [63:0] matmult_in_a71,
    input wire signed [63:0] matmult_in_a72,
    input wire signed [63:0] matmult_in_a73,
    input wire signed [63:0] matmult_in_a74,
    input wire signed [63:0] matmult_in_a75,
    input wire signed [63:0] matmult_in_a76,
    input wire signed [63:0] matmult_in_a77,
    input wire signed [63:0] matmult_in_a78,
    input wire signed [63:0] matmult_in_a79,
    input wire signed [63:0] matmult_in_a80,
    input wire signed [63:0] matmult_in_a81,
    input wire signed [63:0] matmult_in_a82,
    input wire signed [63:0] matmult_in_a83,
    input wire signed [63:0] matmult_in_a84,
    input wire signed [63:0] matmult_in_a85,
    input wire signed [63:0] matmult_in_a86,
    input wire signed [63:0] matmult_in_a87,
    input wire signed [63:0] matmult_in_a88,
    input wire signed [63:0] matmult_in_a89,
    input wire signed [63:0] matmult_in_a90,
    input wire signed [63:0] matmult_in_a91,
    input wire signed [63:0] matmult_in_a92,
    input wire signed [63:0] matmult_in_a93,
    input wire signed [63:0] matmult_in_a94,
    input wire signed [63:0] matmult_in_a95,
    input wire signed [63:0] matmult_in_a96,
    input wire signed [63:0] matmult_in_a97,
    input wire signed [63:0] matmult_in_a98,
    input wire signed [63:0] matmult_in_a99,
    input wire signed [63:0] matmult_in_a100,
    input wire signed [63:0] matmult_in_a101,
    input wire signed [63:0] matmult_in_a102,
    input wire signed [63:0] matmult_in_a103,
    input wire signed [63:0] matmult_in_a104,
    input wire signed [63:0] matmult_in_a105,
    input wire signed [63:0] matmult_in_a106,
    input wire signed [63:0] matmult_in_a107,
    input wire signed [63:0] matmult_in_a108,
    input wire signed [63:0] matmult_in_a109,
    input wire signed [63:0] matmult_in_a110,
    input wire signed [63:0] matmult_in_a111,
    input wire signed [63:0] matmult_in_a112,
    input wire signed [63:0] matmult_in_a113,
    input wire signed [63:0] matmult_in_a114,
    input wire signed [63:0] matmult_in_a115,
    input wire signed [63:0] matmult_in_a116,
    input wire signed [63:0] matmult_in_a117,
    input wire signed [63:0] matmult_in_a118,
    input wire signed [63:0] matmult_in_a119,
    input wire signed [63:0] matmult_in_a120,
    input wire signed [63:0] matmult_in_a121,
    input wire signed [63:0] matmult_in_a122,
    input wire signed [63:0] matmult_in_a123,
    input wire signed [63:0] matmult_in_a124,
    input wire signed [63:0] matmult_in_a125,
    input wire signed [63:0] matmult_in_a126,
    input wire signed [63:0] matmult_in_a127,
    input wire signed [63:0] matmult_in_a128,
    input wire signed [63:0] matmult_in_a129,
    input wire signed [63:0] matmult_in_a130,
    input wire signed [63:0] matmult_in_a131,
    input wire signed [63:0] matmult_in_a132,
    input wire signed [63:0] matmult_in_a133,
    input wire signed [63:0] matmult_in_a134,
    input wire signed [63:0] matmult_in_a135,
    input wire signed [63:0] matmult_in_a136,
    input wire signed [63:0] matmult_in_a137,
    input wire signed [63:0] matmult_in_a138,
    input wire signed [63:0] matmult_in_a139,
    input wire signed [63:0] matmult_in_a140,
    input wire signed [63:0] matmult_in_a141,
    input wire signed [63:0] matmult_in_a142,
    input wire signed [63:0] matmult_in_a143,
    input wire signed [63:0] matmult_in_a144,
    input wire signed [63:0] matmult_in_a145,
    input wire signed [63:0] matmult_in_a146,
    input wire signed [63:0] matmult_in_a147,
    input wire signed [63:0] matmult_in_a148,
    input wire signed [63:0] matmult_in_a149,
    input wire signed [63:0] matmult_in_a150,
    input wire signed [63:0] matmult_in_a151,
    input wire signed [63:0] matmult_in_a152,
    input wire signed [63:0] matmult_in_a153,
    input wire signed [63:0] matmult_in_a154,
    input wire signed [63:0] matmult_in_a155,
    input wire signed [63:0] matmult_in_a156,
    input wire signed [63:0] matmult_in_a157,
    input wire signed [63:0] matmult_in_a158,
    input wire signed [63:0] matmult_in_a159,
    input wire signed [63:0] matmult_in_a160,
    input wire signed [63:0] matmult_in_a161,
    input wire signed [63:0] matmult_in_a162,
    input wire signed [63:0] matmult_in_a163,
    input wire signed [63:0] matmult_in_a164,
    input wire signed [63:0] matmult_in_a165,
    input wire signed [63:0] matmult_in_a166,
    input wire signed [63:0] matmult_in_a167,
    input wire signed [63:0] matmult_in_a168,
    input wire signed [63:0] matmult_in_a169,
    input wire signed [63:0] matmult_in_a170,
    input wire signed [63:0] matmult_in_a171,
    input wire signed [63:0] matmult_in_a172,
    input wire signed [63:0] matmult_in_a173,
    input wire signed [63:0] matmult_in_a174,
    input wire signed [63:0] matmult_in_a175,
    input wire signed [63:0] matmult_in_a176,
    input wire signed [63:0] matmult_in_a177,
    input wire signed [63:0] matmult_in_a178,
    input wire signed [63:0] matmult_in_a179,
    input wire signed [63:0] matmult_in_a180,
    input wire signed [63:0] matmult_in_a181,
    input wire signed [63:0] matmult_in_a182,
    input wire signed [63:0] matmult_in_a183,
    input wire signed [63:0] matmult_in_a184,
    input wire signed [63:0] matmult_in_a185,
    input wire signed [63:0] matmult_in_a186,
    input wire signed [63:0] matmult_in_a187,
    input wire signed [63:0] matmult_in_a188,
    input wire signed [63:0] matmult_in_a189,
    input wire signed [63:0] matmult_in_a190,
    input wire signed [63:0] matmult_in_a191,
    input wire signed [63:0] matmult_in_a192,
    input wire signed [63:0] matmult_in_a193,
    input wire signed [63:0] matmult_in_a194,
    input wire signed [63:0] matmult_in_a195,
    input wire signed [63:0] matmult_in_a196,
    input wire signed [63:0] matmult_in_a197,
    input wire signed [63:0] matmult_in_a198,
    input wire signed [63:0] matmult_in_a199,
    input wire signed [63:0] matmult_in_a200,
    input wire signed [63:0] matmult_in_a201,
    input wire signed [63:0] matmult_in_a202,
    input wire signed [63:0] matmult_in_a203,
    input wire signed [63:0] matmult_in_a204,
    input wire signed [63:0] matmult_in_a205,
    input wire signed [63:0] matmult_in_a206,
    input wire signed [63:0] matmult_in_a207,
    input wire signed [63:0] matmult_in_a208,
    input wire signed [63:0] matmult_in_a209,
    input wire signed [63:0] matmult_in_a210,
    input wire signed [63:0] matmult_in_a211,
    input wire signed [63:0] matmult_in_a212,
    input wire signed [63:0] matmult_in_a213,
    input wire signed [63:0] matmult_in_a214,
    input wire signed [63:0] matmult_in_a215,
    input wire signed [63:0] matmult_in_a216,
    input wire signed [63:0] matmult_in_a217,
    input wire signed [63:0] matmult_in_a218,
    input wire signed [63:0] matmult_in_a219,
    input wire signed [63:0] matmult_in_a220,
    input wire signed [63:0] matmult_in_a221,
    input wire signed [63:0] matmult_in_a222,
    input wire signed [63:0] matmult_in_a223,
    input wire signed [63:0] matmult_in_a224,
    input wire signed [63:0] matmult_in_a225,
    input wire signed [63:0] matmult_in_a226,
    input wire signed [63:0] matmult_in_a227,
    input wire signed [63:0] matmult_in_a228,
    input wire signed [63:0] matmult_in_a229,
    input wire signed [63:0] matmult_in_a230,
    input wire signed [63:0] matmult_in_a231,
    input wire signed [63:0] matmult_in_a232,
    input wire signed [63:0] matmult_in_a233,
    input wire signed [63:0] matmult_in_a234,
    input wire signed [63:0] matmult_in_a235,
    input wire signed [63:0] matmult_in_a236,
    input wire signed [63:0] matmult_in_a237,
    input wire signed [63:0] matmult_in_a238,
    input wire signed [63:0] matmult_in_a239,
    input wire signed [63:0] matmult_in_a240,
    input wire signed [63:0] matmult_in_a241,
    input wire signed [63:0] matmult_in_a242,
    input wire signed [63:0] matmult_in_a243,
    input wire signed [63:0] matmult_in_a244,
    input wire signed [63:0] matmult_in_a245,
    input wire signed [63:0] matmult_in_a246,
    input wire signed [63:0] matmult_in_a247,
    input wire signed [63:0] matmult_in_a248,
    input wire signed [63:0] matmult_in_a249,
    input wire signed [63:0] matmult_in_a250,
    input wire signed [63:0] matmult_in_a251,
    input wire signed [63:0] matmult_in_a252,
    input wire signed [63:0] matmult_in_a253,
    input wire signed [63:0] matmult_in_a254,
    input wire signed [63:0] matmult_in_a255,
    input wire signed [63:0] matmult_in_a256,
    input wire signed [63:0] matmult_in_a257,
    input wire signed [63:0] matmult_in_a258,
    input wire signed [63:0] matmult_in_a259,
    input wire signed [63:0] matmult_in_a260,
    input wire signed [63:0] matmult_in_a261,
    input wire signed [63:0] matmult_in_a262,
    input wire signed [63:0] matmult_in_a263,
    input wire signed [63:0] matmult_in_a264,
    input wire signed [63:0] matmult_in_a265,
    input wire signed [63:0] matmult_in_a266,
    input wire signed [63:0] matmult_in_a267,
    input wire signed [63:0] matmult_in_a268,
    input wire signed [63:0] matmult_in_a269,
    input wire signed [63:0] matmult_in_a270,
    input wire signed [63:0] matmult_in_a271,
    input wire signed [63:0] matmult_in_a272,
    input wire signed [63:0] matmult_in_a273,
    input wire signed [63:0] matmult_in_a274,
    input wire signed [63:0] matmult_in_a275,
    input wire signed [63:0] matmult_in_a276,
    input wire signed [63:0] matmult_in_a277,
    input wire signed [63:0] matmult_in_a278,
    input wire signed [63:0] matmult_in_a279,
    output wire signed [63:0] matmult_out_a0,
    output wire signed [63:0] matmult_out_a1,
    output wire signed [63:0] matmult_out_a2,
    output wire signed [63:0] matmult_out_a3,
    output wire signed [63:0] matmult_out_a4,
    output wire signed [63:0] matmult_out_a5,
    output wire signed [63:0] matmult_out_a6,
    output wire signed [63:0] matmult_out_a7,
    output wire signed [63:0] matmult_out_a8,
    output wire signed [63:0] matmult_out_a9,
    output wire signed [63:0] matmult_out_a10,
    output wire signed [63:0] matmult_out_a11,
    output wire signed [63:0] matmult_out_a12,
    output wire signed [63:0] matmult_out_a13,
    output wire signed [63:0] matmult_out_a14,
    output wire signed [63:0] matmult_out_a15,
    output wire signed [63:0] matmult_out_a16,
    output wire signed [63:0] matmult_out_a17,
    output wire signed [63:0] matmult_out_a18,
    output wire signed [63:0] matmult_out_a19,
    output wire signed [63:0] matmult_out_a20,
    output wire signed [63:0] matmult_out_a21,
    output wire signed [63:0] matmult_out_a22,
    output wire signed [63:0] matmult_out_a23,
    output wire signed [63:0] matmult_out_a24,
    output wire signed [63:0] matmult_out_a25,
    output wire signed [63:0] matmult_out_a26,
    output wire signed [63:0] matmult_out_a27,
    output wire signed [63:0] matmult_out_a28,
    output wire signed [63:0] matmult_out_a29,
    output wire signed [63:0] matmult_out_a30,
    output wire signed [63:0] matmult_out_a31,
    output wire signed [63:0] matmult_out_a32,
    output wire signed [63:0] matmult_out_a33,
    output wire signed [63:0] matmult_out_a34,
    output wire signed [63:0] matmult_out_a35,
    output wire signed [63:0] matmult_out_a36,
    output wire signed [63:0] matmult_out_a37,
    output wire signed [63:0] matmult_out_a38,
    output wire signed [63:0] matmult_out_a39,
    output wire signed [63:0] matmult_out_a40,
    output wire signed [63:0] matmult_out_a41,
    output wire signed [63:0] matmult_out_a42,
    output wire signed [63:0] matmult_out_a43,
    output wire signed [63:0] matmult_out_a44,
    output wire signed [63:0] matmult_out_a45,
    output wire signed [63:0] matmult_out_a46,
    output wire signed [63:0] matmult_out_a47,
    output wire signed [63:0] matmult_out_a48,
    output wire signed [63:0] matmult_out_a49,
    output wire signed [63:0] matmult_out_a50,
    output wire signed [63:0] matmult_out_a51,
    output wire signed [63:0] matmult_out_a52,
    output wire signed [63:0] matmult_out_a53,
    output wire signed [63:0] matmult_out_a54,
    output wire signed [63:0] matmult_out_a55,
    output wire signed [63:0] matmult_out_a56,
    output wire signed [63:0] matmult_out_a57,
    output wire signed [63:0] matmult_out_a58,
    output wire signed [63:0] matmult_out_a59,
    output wire signed [63:0] matmult_out_a60,
    output wire signed [63:0] matmult_out_a61,
    output wire signed [63:0] matmult_out_a62,
    output wire signed [63:0] matmult_out_a63,
    output wire signed [63:0] matmult_out_a64,
    output wire signed [63:0] matmult_out_a65,
    output wire signed [63:0] matmult_out_a66,
    output wire signed [63:0] matmult_out_a67,
    output wire signed [63:0] matmult_out_a68,
    output wire signed [63:0] matmult_out_a69,
    output wire signed [63:0] matmult_out_a70,
    output wire signed [63:0] matmult_out_a71,
    output wire signed [63:0] matmult_out_a72,
    output wire signed [63:0] matmult_out_a73,
    output wire signed [63:0] matmult_out_a74,
    output wire signed [63:0] matmult_out_a75,
    output wire signed [63:0] matmult_out_a76,
    output wire signed [63:0] matmult_out_a77,
    output wire signed [63:0] matmult_out_a78,
    output wire signed [63:0] matmult_out_a79,
    output wire signed [63:0] matmult_out_a80,
    output wire signed [63:0] matmult_out_a81,
    output wire signed [63:0] matmult_out_a82,
    output wire signed [63:0] matmult_out_a83,
    output wire signed [63:0] matmult_out_a84,
    output wire signed [63:0] matmult_out_a85,
    output wire signed [63:0] matmult_out_a86,
    output wire signed [63:0] matmult_out_a87,
    output wire signed [63:0] matmult_out_a88,
    output wire signed [63:0] matmult_out_a89,
    output wire signed [63:0] matmult_out_a90,
    output wire signed [63:0] matmult_out_a91,
    output wire signed [63:0] matmult_out_a92,
    output wire signed [63:0] matmult_out_a93,
    output wire signed [63:0] matmult_out_a94,
    output wire signed [63:0] matmult_out_a95,
    output wire signed [63:0] matmult_out_a96,
    output wire signed [63:0] matmult_out_a97,
    output wire signed [63:0] matmult_out_a98,
    output wire signed [63:0] matmult_out_a99,
    output wire signed [63:0] matmult_out_a100,
    output wire signed [63:0] matmult_out_a101,
    output wire signed [63:0] matmult_out_a102,
    output wire signed [63:0] matmult_out_a103,
    output wire signed [63:0] matmult_out_a104,
    output wire signed [63:0] matmult_out_a105,
    output wire signed [63:0] matmult_out_a106,
    output wire signed [63:0] matmult_out_a107,
    output wire signed [63:0] matmult_out_a108,
    output wire signed [63:0] matmult_out_a109,
    output wire signed [63:0] matmult_out_a110,
    output wire signed [63:0] matmult_out_a111,
    output wire signed [63:0] matmult_out_a112,
    output wire signed [63:0] matmult_out_a113,
    output wire signed [63:0] matmult_out_a114,
    output wire signed [63:0] matmult_out_a115,
    output wire signed [63:0] matmult_out_a116,
    output wire signed [63:0] matmult_out_a117,
    output wire signed [63:0] matmult_out_a118,
    output wire signed [63:0] matmult_out_a119,
    output wire signed [63:0] matmult_out_a120,
    output wire signed [63:0] matmult_out_a121,
    output wire signed [63:0] matmult_out_a122,
    output wire signed [63:0] matmult_out_a123,
    output wire signed [63:0] matmult_out_a124,
    output wire signed [63:0] matmult_out_a125,
    output wire signed [63:0] matmult_out_a126,
    output wire signed [63:0] matmult_out_a127,
    output wire signed [63:0] matmult_out_a128,
    output wire signed [63:0] matmult_out_a129,
    output wire signed [63:0] matmult_out_a130,
    output wire signed [63:0] matmult_out_a131,
    output wire signed [63:0] matmult_out_a132,
    output wire signed [63:0] matmult_out_a133,
    output wire signed [63:0] matmult_out_a134,
    output wire signed [63:0] matmult_out_a135,
    output wire signed [63:0] matmult_out_a136,
    output wire signed [63:0] matmult_out_a137,
    output wire signed [63:0] matmult_out_a138,
    output wire signed [63:0] matmult_out_a139,
    output wire signed [63:0] matmult_out_a140,
    output wire signed [63:0] matmult_out_a141,
    output wire signed [63:0] matmult_out_a142,
    output wire signed [63:0] matmult_out_a143,
    output wire signed [63:0] matmult_out_a144,
    output wire signed [63:0] matmult_out_a145,
    output wire signed [63:0] matmult_out_a146,
    output wire signed [63:0] matmult_out_a147,
    output wire signed [63:0] matmult_out_a148,
    output wire signed [63:0] matmult_out_a149,
    output wire signed [63:0] matmult_out_a150,
    output wire signed [63:0] matmult_out_a151,
    output wire signed [63:0] matmult_out_a152,
    output wire signed [63:0] matmult_out_a153,
    output wire signed [63:0] matmult_out_a154,
    output wire signed [63:0] matmult_out_a155,
    output wire signed [63:0] matmult_out_a156,
    output wire signed [63:0] matmult_out_a157,
    output wire signed [63:0] matmult_out_a158,
    output wire signed [63:0] matmult_out_a159,
    output wire signed [63:0] matmult_out_a160,
    output wire signed [63:0] matmult_out_a161,
    output wire signed [63:0] matmult_out_a162,
    output wire signed [63:0] matmult_out_a163,
    output wire signed [63:0] matmult_out_a164,
    output wire signed [63:0] matmult_out_a165,
    output wire signed [63:0] matmult_out_a166,
    output wire signed [63:0] matmult_out_a167,
    output wire signed [63:0] matmult_out_a168,
    output wire signed [63:0] matmult_out_a169,
    output wire signed [63:0] matmult_out_a170,
    output wire signed [63:0] matmult_out_a171,
    output wire signed [63:0] matmult_out_a172,
    output wire signed [63:0] matmult_out_a173,
    output wire signed [63:0] matmult_out_a174,
    output wire signed [63:0] matmult_out_a175,
    output wire signed [63:0] matmult_out_a176,
    output wire signed [63:0] matmult_out_a177,
    output wire signed [63:0] matmult_out_a178,
    output wire signed [63:0] matmult_out_a179,
    output wire signed [63:0] matmult_out_a180,
    output wire signed [63:0] matmult_out_a181,
    output wire signed [63:0] matmult_out_a182,
    output wire signed [63:0] matmult_out_a183,
    output wire signed [63:0] matmult_out_a184,
    output wire signed [63:0] matmult_out_a185,
    output wire signed [63:0] matmult_out_a186,
    output wire signed [63:0] matmult_out_a187,
    output wire signed [63:0] matmult_out_a188,
    output wire signed [63:0] matmult_out_a189,
    output wire signed [63:0] matmult_out_a190,
    output wire signed [63:0] matmult_out_a191,
    output wire signed [63:0] matmult_out_a192,
    output wire signed [63:0] matmult_out_a193,
    output wire signed [63:0] matmult_out_a194,
    output wire signed [63:0] matmult_out_a195,
    output wire signed [63:0] matmult_out_a196,
    output wire signed [63:0] matmult_out_a197,
    output wire signed [63:0] matmult_out_a198,
    output wire signed [63:0] matmult_out_a199,
    output wire signed [63:0] matmult_out_a200,
    output wire signed [63:0] matmult_out_a201,
    output wire signed [63:0] matmult_out_a202,
    output wire signed [63:0] matmult_out_a203,
    output wire signed [63:0] matmult_out_a204,
    output wire signed [63:0] matmult_out_a205,
    output wire signed [63:0] matmult_out_a206,
    output wire signed [63:0] matmult_out_a207,
    output wire signed [63:0] matmult_out_a208,
    output wire signed [63:0] matmult_out_a209,
    output wire signed [63:0] matmult_out_a210,
    output wire signed [63:0] matmult_out_a211,
    output wire signed [63:0] matmult_out_a212,
    output wire signed [63:0] matmult_out_a213,
    output wire signed [63:0] matmult_out_a214,
    output wire signed [63:0] matmult_out_a215,
    output wire signed [63:0] matmult_out_a216,
    output wire signed [63:0] matmult_out_a217,
    output wire signed [63:0] matmult_out_a218,
    output wire signed [63:0] matmult_out_a219,
    output wire signed [63:0] matmult_out_a220,
    output wire signed [63:0] matmult_out_a221,
    output wire signed [63:0] matmult_out_a222,
    output wire signed [63:0] matmult_out_a223,
    output wire signed [63:0] matmult_out_a224,
    output wire signed [63:0] matmult_out_a225,
    output wire signed [63:0] matmult_out_a226,
    output wire signed [63:0] matmult_out_a227,
    output wire signed [63:0] matmult_out_a228,
    output wire signed [63:0] matmult_out_a229,
    output wire signed [63:0] matmult_out_a230,
    output wire signed [63:0] matmult_out_a231,
    output wire signed [63:0] matmult_out_a232,
    output wire signed [63:0] matmult_out_a233,
    output wire signed [63:0] matmult_out_a234,
    output wire signed [63:0] matmult_out_a235,
    output wire signed [63:0] matmult_out_a236,
    output wire signed [63:0] matmult_out_a237,
    output wire signed [63:0] matmult_out_a238,
    output wire signed [63:0] matmult_out_a239,
    output wire signed [63:0] matmult_out_a240,
    output wire signed [63:0] matmult_out_a241,
    output wire signed [63:0] matmult_out_a242,
    output wire signed [63:0] matmult_out_a243,
    output wire signed [63:0] matmult_out_a244,
    output wire signed [63:0] matmult_out_a245,
    output wire signed [63:0] matmult_out_a246,
    output wire signed [63:0] matmult_out_a247,
    output wire signed [63:0] matmult_out_a248,
    output wire signed [63:0] matmult_out_a249,
    output wire signed [63:0] matmult_out_a250,
    output wire signed [63:0] matmult_out_a251,
    output wire signed [63:0] matmult_out_a252,
    output wire signed [63:0] matmult_out_a253,
    output wire signed [63:0] matmult_out_a254,
    output wire signed [63:0] matmult_out_a255,
    output wire signed [63:0] matmult_out_a256,
    output wire signed [63:0] matmult_out_a257,
    output wire signed [63:0] matmult_out_a258,
    output wire signed [63:0] matmult_out_a259,
    output wire signed [63:0] matmult_out_a260,
    output wire signed [63:0] matmult_out_a261,
    output wire signed [63:0] matmult_out_a262,
    output wire signed [63:0] matmult_out_a263,
    output wire signed [63:0] matmult_out_a264,
    output wire signed [63:0] matmult_out_a265,
    output wire signed [63:0] matmult_out_a266,
    output wire signed [63:0] matmult_out_a267,
    output wire signed [63:0] matmult_out_a268,
    output wire signed [63:0] matmult_out_a269,
    output wire signed [63:0] matmult_out_a270,
    output wire signed [63:0] matmult_out_a271,
    output wire signed [63:0] matmult_out_a272,
    output wire signed [63:0] matmult_out_a273,
    output wire signed [63:0] matmult_out_a274,
    output wire signed [63:0] matmult_out_a275,
    output wire signed [63:0] matmult_out_a276,
    output wire signed [63:0] matmult_out_a277,
    output wire signed [63:0] matmult_out_a278,
    output wire signed [63:0] matmult_out_a279,
    input wire signed [63:0] matmult_in_b0,
    input wire signed [63:0] matmult_in_b1,
    input wire signed [63:0] matmult_in_b2,
    input wire signed [63:0] matmult_in_b3,
    input wire signed [63:0] matmult_in_b4,
    input wire signed [63:0] matmult_in_b5,
    input wire signed [63:0] matmult_in_b6,
    input wire signed [63:0] matmult_in_b7,
    input wire signed [63:0] matmult_in_b8,
    input wire signed [63:0] matmult_in_b9,
    input wire signed [63:0] matmult_in_b10,
    input wire signed [63:0] matmult_in_b11,
    input wire signed [63:0] matmult_in_b12,
    input wire signed [63:0] matmult_in_b13,
    input wire signed [63:0] matmult_in_b14,
    input wire signed [63:0] matmult_in_b15,
    input wire signed [63:0] matmult_in_b16,
    input wire signed [63:0] matmult_in_b17,
    input wire signed [63:0] matmult_in_b18,
    input wire signed [63:0] matmult_in_b19,
    input wire signed [63:0] matmult_in_b20,
    input wire signed [63:0] matmult_in_b21,
    input wire signed [63:0] matmult_in_b22,
    input wire signed [63:0] matmult_in_b23,
    input wire signed [63:0] matmult_in_b24,
    input wire signed [63:0] matmult_in_b25,
    input wire signed [63:0] matmult_in_b26,
    input wire signed [63:0] matmult_in_b27,
    input wire signed [63:0] matmult_in_b28,
    input wire signed [63:0] matmult_in_b29,
    input wire signed [63:0] matmult_in_b30,
    input wire signed [63:0] matmult_in_b31,
    input wire signed [63:0] matmult_in_b32,
    input wire signed [63:0] matmult_in_b33,
    input wire signed [63:0] matmult_in_b34,
    input wire signed [63:0] matmult_in_b35,
    input wire signed [63:0] matmult_in_b36,
    input wire signed [63:0] matmult_in_b37,
    input wire signed [63:0] matmult_in_b38,
    input wire signed [63:0] matmult_in_b39,
    input wire signed [63:0] matmult_in_b40,
    input wire signed [63:0] matmult_in_b41,
    input wire signed [63:0] matmult_in_b42,
    input wire signed [63:0] matmult_in_b43,
    input wire signed [63:0] matmult_in_b44,
    input wire signed [63:0] matmult_in_b45,
    input wire signed [63:0] matmult_in_b46,
    input wire signed [63:0] matmult_in_b47,
    input wire signed [63:0] matmult_in_b48,
    input wire signed [63:0] matmult_in_b49,
    input wire signed [63:0] matmult_in_b50,
    input wire signed [63:0] matmult_in_b51,
    input wire signed [63:0] matmult_in_b52,
    input wire signed [63:0] matmult_in_b53,
    input wire signed [63:0] matmult_in_b54,
    input wire signed [63:0] matmult_in_b55,
    input wire signed [63:0] matmult_in_b56,
    input wire signed [63:0] matmult_in_b57,
    input wire signed [63:0] matmult_in_b58,
    input wire signed [63:0] matmult_in_b59,
    input wire signed [63:0] matmult_in_b60,
    input wire signed [63:0] matmult_in_b61,
    input wire signed [63:0] matmult_in_b62,
    input wire signed [63:0] matmult_in_b63,
    input wire signed [63:0] matmult_in_b64,
    input wire signed [63:0] matmult_in_b65,
    input wire signed [63:0] matmult_in_b66,
    input wire signed [63:0] matmult_in_b67,
    input wire signed [63:0] matmult_in_b68,
    input wire signed [63:0] matmult_in_b69,
    input wire signed [63:0] matmult_in_b70,
    input wire signed [63:0] matmult_in_b71,
    input wire signed [63:0] matmult_in_b72,
    input wire signed [63:0] matmult_in_b73,
    input wire signed [63:0] matmult_in_b74,
    input wire signed [63:0] matmult_in_b75,
    input wire signed [63:0] matmult_in_b76,
    input wire signed [63:0] matmult_in_b77,
    input wire signed [63:0] matmult_in_b78,
    input wire signed [63:0] matmult_in_b79,
    input wire signed [63:0] matmult_in_b80,
    input wire signed [63:0] matmult_in_b81,
    input wire signed [63:0] matmult_in_b82,
    input wire signed [63:0] matmult_in_b83,
    input wire signed [63:0] matmult_in_b84,
    input wire signed [63:0] matmult_in_b85,
    input wire signed [63:0] matmult_in_b86,
    input wire signed [63:0] matmult_in_b87,
    input wire signed [63:0] matmult_in_b88,
    input wire signed [63:0] matmult_in_b89,
    input wire signed [63:0] matmult_in_b90,
    input wire signed [63:0] matmult_in_b91,
    input wire signed [63:0] matmult_in_b92,
    input wire signed [63:0] matmult_in_b93,
    input wire signed [63:0] matmult_in_b94,
    input wire signed [63:0] matmult_in_b95,
    input wire signed [63:0] matmult_in_b96,
    input wire signed [63:0] matmult_in_b97,
    input wire signed [63:0] matmult_in_b98,
    input wire signed [63:0] matmult_in_b99,
    input wire signed [63:0] matmult_in_b100,
    input wire signed [63:0] matmult_in_b101,
    input wire signed [63:0] matmult_in_b102,
    input wire signed [63:0] matmult_in_b103,
    input wire signed [63:0] matmult_in_b104,
    input wire signed [63:0] matmult_in_b105,
    input wire signed [63:0] matmult_in_b106,
    input wire signed [63:0] matmult_in_b107,
    input wire signed [63:0] matmult_in_b108,
    input wire signed [63:0] matmult_in_b109,
    input wire signed [63:0] matmult_in_b110,
    input wire signed [63:0] matmult_in_b111,
    input wire signed [63:0] matmult_in_b112,
    input wire signed [63:0] matmult_in_b113,
    input wire signed [63:0] matmult_in_b114,
    input wire signed [63:0] matmult_in_b115,
    input wire signed [63:0] matmult_in_b116,
    input wire signed [63:0] matmult_in_b117,
    input wire signed [63:0] matmult_in_b118,
    input wire signed [63:0] matmult_in_b119,
    input wire signed [63:0] matmult_in_b120,
    input wire signed [63:0] matmult_in_b121,
    input wire signed [63:0] matmult_in_b122,
    input wire signed [63:0] matmult_in_b123,
    input wire signed [63:0] matmult_in_b124,
    input wire signed [63:0] matmult_in_b125,
    input wire signed [63:0] matmult_in_b126,
    input wire signed [63:0] matmult_in_b127,
    input wire signed [63:0] matmult_in_b128,
    input wire signed [63:0] matmult_in_b129,
    input wire signed [63:0] matmult_in_b130,
    input wire signed [63:0] matmult_in_b131,
    input wire signed [63:0] matmult_in_b132,
    input wire signed [63:0] matmult_in_b133,
    input wire signed [63:0] matmult_in_b134,
    input wire signed [63:0] matmult_in_b135,
    input wire signed [63:0] matmult_in_b136,
    input wire signed [63:0] matmult_in_b137,
    input wire signed [63:0] matmult_in_b138,
    input wire signed [63:0] matmult_in_b139,
    input wire signed [63:0] matmult_in_b140,
    input wire signed [63:0] matmult_in_b141,
    input wire signed [63:0] matmult_in_b142,
    input wire signed [63:0] matmult_in_b143,
    input wire signed [63:0] matmult_in_b144,
    input wire signed [63:0] matmult_in_b145,
    input wire signed [63:0] matmult_in_b146,
    input wire signed [63:0] matmult_in_b147,
    input wire signed [63:0] matmult_in_b148,
    input wire signed [63:0] matmult_in_b149,
    input wire signed [63:0] matmult_in_b150,
    input wire signed [63:0] matmult_in_b151,
    input wire signed [63:0] matmult_in_b152,
    input wire signed [63:0] matmult_in_b153,
    input wire signed [63:0] matmult_in_b154,
    input wire signed [63:0] matmult_in_b155,
    input wire signed [63:0] matmult_in_b156,
    input wire signed [63:0] matmult_in_b157,
    input wire signed [63:0] matmult_in_b158,
    input wire signed [63:0] matmult_in_b159,
    input wire signed [63:0] matmult_in_b160,
    input wire signed [63:0] matmult_in_b161,
    input wire signed [63:0] matmult_in_b162,
    input wire signed [63:0] matmult_in_b163,
    input wire signed [63:0] matmult_in_b164,
    input wire signed [63:0] matmult_in_b165,
    input wire signed [63:0] matmult_in_b166,
    input wire signed [63:0] matmult_in_b167,
    input wire signed [63:0] matmult_in_b168,
    input wire signed [63:0] matmult_in_b169,
    input wire signed [63:0] matmult_in_b170,
    input wire signed [63:0] matmult_in_b171,
    input wire signed [63:0] matmult_in_b172,
    input wire signed [63:0] matmult_in_b173,
    input wire signed [63:0] matmult_in_b174,
    input wire signed [63:0] matmult_in_b175,
    input wire signed [63:0] matmult_in_b176,
    input wire signed [63:0] matmult_in_b177,
    input wire signed [63:0] matmult_in_b178,
    input wire signed [63:0] matmult_in_b179,
    input wire signed [63:0] matmult_in_b180,
    input wire signed [63:0] matmult_in_b181,
    input wire signed [63:0] matmult_in_b182,
    input wire signed [63:0] matmult_in_b183,
    input wire signed [63:0] matmult_in_b184,
    input wire signed [63:0] matmult_in_b185,
    input wire signed [63:0] matmult_in_b186,
    input wire signed [63:0] matmult_in_b187,
    input wire signed [63:0] matmult_in_b188,
    input wire signed [63:0] matmult_in_b189,
    input wire signed [63:0] matmult_in_b190,
    input wire signed [63:0] matmult_in_b191,
    input wire signed [63:0] matmult_in_b192,
    input wire signed [63:0] matmult_in_b193,
    input wire signed [63:0] matmult_in_b194,
    input wire signed [63:0] matmult_in_b195,
    input wire signed [63:0] matmult_in_b196,
    input wire signed [63:0] matmult_in_b197,
    input wire signed [63:0] matmult_in_b198,
    input wire signed [63:0] matmult_in_b199,
    input wire signed [63:0] matmult_in_b200,
    input wire signed [63:0] matmult_in_b201,
    input wire signed [63:0] matmult_in_b202,
    input wire signed [63:0] matmult_in_b203,
    input wire signed [63:0] matmult_in_b204,
    input wire signed [63:0] matmult_in_b205,
    input wire signed [63:0] matmult_in_b206,
    input wire signed [63:0] matmult_in_b207,
    input wire signed [63:0] matmult_in_b208,
    input wire signed [63:0] matmult_in_b209,
    input wire signed [63:0] matmult_in_b210,
    input wire signed [63:0] matmult_in_b211,
    input wire signed [63:0] matmult_in_b212,
    input wire signed [63:0] matmult_in_b213,
    input wire signed [63:0] matmult_in_b214,
    input wire signed [63:0] matmult_in_b215,
    input wire signed [63:0] matmult_in_b216,
    input wire signed [63:0] matmult_in_b217,
    input wire signed [63:0] matmult_in_b218,
    input wire signed [63:0] matmult_in_b219,
    input wire signed [63:0] matmult_in_b220,
    input wire signed [63:0] matmult_in_b221,
    input wire signed [63:0] matmult_in_b222,
    input wire signed [63:0] matmult_in_b223,
    input wire signed [63:0] matmult_in_b224,
    input wire signed [63:0] matmult_in_b225,
    input wire signed [63:0] matmult_in_b226,
    input wire signed [63:0] matmult_in_b227,
    input wire signed [63:0] matmult_in_b228,
    input wire signed [63:0] matmult_in_b229,
    input wire signed [63:0] matmult_in_b230,
    input wire signed [63:0] matmult_in_b231,
    input wire signed [63:0] matmult_in_b232,
    input wire signed [63:0] matmult_in_b233,
    input wire signed [63:0] matmult_in_b234,
    input wire signed [63:0] matmult_in_b235,
    input wire signed [63:0] matmult_in_b236,
    input wire signed [63:0] matmult_in_b237,
    input wire signed [63:0] matmult_in_b238,
    input wire signed [63:0] matmult_in_b239,
    input wire signed [63:0] matmult_in_b240,
    input wire signed [63:0] matmult_in_b241,
    input wire signed [63:0] matmult_in_b242,
    input wire signed [63:0] matmult_in_b243,
    input wire signed [63:0] matmult_in_b244,
    input wire signed [63:0] matmult_in_b245,
    input wire signed [63:0] matmult_in_b246,
    input wire signed [63:0] matmult_in_b247,
    input wire signed [63:0] matmult_in_b248,
    input wire signed [63:0] matmult_in_b249,
    input wire signed [63:0] matmult_in_b250,
    input wire signed [63:0] matmult_in_b251,
    input wire signed [63:0] matmult_in_b252,
    input wire signed [63:0] matmult_in_b253,
    input wire signed [63:0] matmult_in_b254,
    input wire signed [63:0] matmult_in_b255,
    input wire signed [63:0] matmult_in_b256,
    input wire signed [63:0] matmult_in_b257,
    input wire signed [63:0] matmult_in_b258,
    input wire signed [63:0] matmult_in_b259,
    input wire signed [63:0] matmult_in_b260,
    input wire signed [63:0] matmult_in_b261,
    input wire signed [63:0] matmult_in_b262,
    input wire signed [63:0] matmult_in_b263,
    input wire signed [63:0] matmult_in_b264,
    input wire signed [63:0] matmult_in_b265,
    input wire signed [63:0] matmult_in_b266,
    input wire signed [63:0] matmult_in_b267,
    input wire signed [63:0] matmult_in_b268,
    input wire signed [63:0] matmult_in_b269,
    input wire signed [63:0] matmult_in_b270,
    input wire signed [63:0] matmult_in_b271,
    input wire signed [63:0] matmult_in_b272,
    input wire signed [63:0] matmult_in_b273,
    input wire signed [63:0] matmult_in_b274,
    input wire signed [63:0] matmult_in_b275,
    input wire signed [63:0] matmult_in_b276,
    input wire signed [63:0] matmult_in_b277,
    input wire signed [63:0] matmult_in_b278,
    input wire signed [63:0] matmult_in_b279,
    output wire signed [63:0] matmult_out_b0,
    output wire signed [63:0] matmult_out_b1,
    output wire signed [63:0] matmult_out_b2,
    output wire signed [63:0] matmult_out_b3,
    output wire signed [63:0] matmult_out_b4,
    output wire signed [63:0] matmult_out_b5,
    output wire signed [63:0] matmult_out_b6,
    output wire signed [63:0] matmult_out_b7,
    output wire signed [63:0] matmult_out_b8,
    output wire signed [63:0] matmult_out_b9,
    output wire signed [63:0] matmult_out_b10,
    output wire signed [63:0] matmult_out_b11,
    output wire signed [63:0] matmult_out_b12,
    output wire signed [63:0] matmult_out_b13,
    output wire signed [63:0] matmult_out_b14,
    output wire signed [63:0] matmult_out_b15,
    output wire signed [63:0] matmult_out_b16,
    output wire signed [63:0] matmult_out_b17,
    output wire signed [63:0] matmult_out_b18,
    output wire signed [63:0] matmult_out_b19,
    output wire signed [63:0] matmult_out_b20,
    output wire signed [63:0] matmult_out_b21,
    output wire signed [63:0] matmult_out_b22,
    output wire signed [63:0] matmult_out_b23,
    output wire signed [63:0] matmult_out_b24,
    output wire signed [63:0] matmult_out_b25,
    output wire signed [63:0] matmult_out_b26,
    output wire signed [63:0] matmult_out_b27,
    output wire signed [63:0] matmult_out_b28,
    output wire signed [63:0] matmult_out_b29,
    output wire signed [63:0] matmult_out_b30,
    output wire signed [63:0] matmult_out_b31,
    output wire signed [63:0] matmult_out_b32,
    output wire signed [63:0] matmult_out_b33,
    output wire signed [63:0] matmult_out_b34,
    output wire signed [63:0] matmult_out_b35,
    output wire signed [63:0] matmult_out_b36,
    output wire signed [63:0] matmult_out_b37,
    output wire signed [63:0] matmult_out_b38,
    output wire signed [63:0] matmult_out_b39,
    output wire signed [63:0] matmult_out_b40,
    output wire signed [63:0] matmult_out_b41,
    output wire signed [63:0] matmult_out_b42,
    output wire signed [63:0] matmult_out_b43,
    output wire signed [63:0] matmult_out_b44,
    output wire signed [63:0] matmult_out_b45,
    output wire signed [63:0] matmult_out_b46,
    output wire signed [63:0] matmult_out_b47,
    output wire signed [63:0] matmult_out_b48,
    output wire signed [63:0] matmult_out_b49,
    output wire signed [63:0] matmult_out_b50,
    output wire signed [63:0] matmult_out_b51,
    output wire signed [63:0] matmult_out_b52,
    output wire signed [63:0] matmult_out_b53,
    output wire signed [63:0] matmult_out_b54,
    output wire signed [63:0] matmult_out_b55,
    output wire signed [63:0] matmult_out_b56,
    output wire signed [63:0] matmult_out_b57,
    output wire signed [63:0] matmult_out_b58,
    output wire signed [63:0] matmult_out_b59,
    output wire signed [63:0] matmult_out_b60,
    output wire signed [63:0] matmult_out_b61,
    output wire signed [63:0] matmult_out_b62,
    output wire signed [63:0] matmult_out_b63,
    output wire signed [63:0] matmult_out_b64,
    output wire signed [63:0] matmult_out_b65,
    output wire signed [63:0] matmult_out_b66,
    output wire signed [63:0] matmult_out_b67,
    output wire signed [63:0] matmult_out_b68,
    output wire signed [63:0] matmult_out_b69,
    output wire signed [63:0] matmult_out_b70,
    output wire signed [63:0] matmult_out_b71,
    output wire signed [63:0] matmult_out_b72,
    output wire signed [63:0] matmult_out_b73,
    output wire signed [63:0] matmult_out_b74,
    output wire signed [63:0] matmult_out_b75,
    output wire signed [63:0] matmult_out_b76,
    output wire signed [63:0] matmult_out_b77,
    output wire signed [63:0] matmult_out_b78,
    output wire signed [63:0] matmult_out_b79,
    output wire signed [63:0] matmult_out_b80,
    output wire signed [63:0] matmult_out_b81,
    output wire signed [63:0] matmult_out_b82,
    output wire signed [63:0] matmult_out_b83,
    output wire signed [63:0] matmult_out_b84,
    output wire signed [63:0] matmult_out_b85,
    output wire signed [63:0] matmult_out_b86,
    output wire signed [63:0] matmult_out_b87,
    output wire signed [63:0] matmult_out_b88,
    output wire signed [63:0] matmult_out_b89,
    output wire signed [63:0] matmult_out_b90,
    output wire signed [63:0] matmult_out_b91,
    output wire signed [63:0] matmult_out_b92,
    output wire signed [63:0] matmult_out_b93,
    output wire signed [63:0] matmult_out_b94,
    output wire signed [63:0] matmult_out_b95,
    output wire signed [63:0] matmult_out_b96,
    output wire signed [63:0] matmult_out_b97,
    output wire signed [63:0] matmult_out_b98,
    output wire signed [63:0] matmult_out_b99,
    output wire signed [63:0] matmult_out_b100,
    output wire signed [63:0] matmult_out_b101,
    output wire signed [63:0] matmult_out_b102,
    output wire signed [63:0] matmult_out_b103,
    output wire signed [63:0] matmult_out_b104,
    output wire signed [63:0] matmult_out_b105,
    output wire signed [63:0] matmult_out_b106,
    output wire signed [63:0] matmult_out_b107,
    output wire signed [63:0] matmult_out_b108,
    output wire signed [63:0] matmult_out_b109,
    output wire signed [63:0] matmult_out_b110,
    output wire signed [63:0] matmult_out_b111,
    output wire signed [63:0] matmult_out_b112,
    output wire signed [63:0] matmult_out_b113,
    output wire signed [63:0] matmult_out_b114,
    output wire signed [63:0] matmult_out_b115,
    output wire signed [63:0] matmult_out_b116,
    output wire signed [63:0] matmult_out_b117,
    output wire signed [63:0] matmult_out_b118,
    output wire signed [63:0] matmult_out_b119,
    output wire signed [63:0] matmult_out_b120,
    output wire signed [63:0] matmult_out_b121,
    output wire signed [63:0] matmult_out_b122,
    output wire signed [63:0] matmult_out_b123,
    output wire signed [63:0] matmult_out_b124,
    output wire signed [63:0] matmult_out_b125,
    output wire signed [63:0] matmult_out_b126,
    output wire signed [63:0] matmult_out_b127,
    output wire signed [63:0] matmult_out_b128,
    output wire signed [63:0] matmult_out_b129,
    output wire signed [63:0] matmult_out_b130,
    output wire signed [63:0] matmult_out_b131,
    output wire signed [63:0] matmult_out_b132,
    output wire signed [63:0] matmult_out_b133,
    output wire signed [63:0] matmult_out_b134,
    output wire signed [63:0] matmult_out_b135,
    output wire signed [63:0] matmult_out_b136,
    output wire signed [63:0] matmult_out_b137,
    output wire signed [63:0] matmult_out_b138,
    output wire signed [63:0] matmult_out_b139,
    output wire signed [63:0] matmult_out_b140,
    output wire signed [63:0] matmult_out_b141,
    output wire signed [63:0] matmult_out_b142,
    output wire signed [63:0] matmult_out_b143,
    output wire signed [63:0] matmult_out_b144,
    output wire signed [63:0] matmult_out_b145,
    output wire signed [63:0] matmult_out_b146,
    output wire signed [63:0] matmult_out_b147,
    output wire signed [63:0] matmult_out_b148,
    output wire signed [63:0] matmult_out_b149,
    output wire signed [63:0] matmult_out_b150,
    output wire signed [63:0] matmult_out_b151,
    output wire signed [63:0] matmult_out_b152,
    output wire signed [63:0] matmult_out_b153,
    output wire signed [63:0] matmult_out_b154,
    output wire signed [63:0] matmult_out_b155,
    output wire signed [63:0] matmult_out_b156,
    output wire signed [63:0] matmult_out_b157,
    output wire signed [63:0] matmult_out_b158,
    output wire signed [63:0] matmult_out_b159,
    output wire signed [63:0] matmult_out_b160,
    output wire signed [63:0] matmult_out_b161,
    output wire signed [63:0] matmult_out_b162,
    output wire signed [63:0] matmult_out_b163,
    output wire signed [63:0] matmult_out_b164,
    output wire signed [63:0] matmult_out_b165,
    output wire signed [63:0] matmult_out_b166,
    output wire signed [63:0] matmult_out_b167,
    output wire signed [63:0] matmult_out_b168,
    output wire signed [63:0] matmult_out_b169,
    output wire signed [63:0] matmult_out_b170,
    output wire signed [63:0] matmult_out_b171,
    output wire signed [63:0] matmult_out_b172,
    output wire signed [63:0] matmult_out_b173,
    output wire signed [63:0] matmult_out_b174,
    output wire signed [63:0] matmult_out_b175,
    output wire signed [63:0] matmult_out_b176,
    output wire signed [63:0] matmult_out_b177,
    output wire signed [63:0] matmult_out_b178,
    output wire signed [63:0] matmult_out_b179,
    output wire signed [63:0] matmult_out_b180,
    output wire signed [63:0] matmult_out_b181,
    output wire signed [63:0] matmult_out_b182,
    output wire signed [63:0] matmult_out_b183,
    output wire signed [63:0] matmult_out_b184,
    output wire signed [63:0] matmult_out_b185,
    output wire signed [63:0] matmult_out_b186,
    output wire signed [63:0] matmult_out_b187,
    output wire signed [63:0] matmult_out_b188,
    output wire signed [63:0] matmult_out_b189,
    output wire signed [63:0] matmult_out_b190,
    output wire signed [63:0] matmult_out_b191,
    output wire signed [63:0] matmult_out_b192,
    output wire signed [63:0] matmult_out_b193,
    output wire signed [63:0] matmult_out_b194,
    output wire signed [63:0] matmult_out_b195,
    output wire signed [63:0] matmult_out_b196,
    output wire signed [63:0] matmult_out_b197,
    output wire signed [63:0] matmult_out_b198,
    output wire signed [63:0] matmult_out_b199,
    output wire signed [63:0] matmult_out_b200,
    output wire signed [63:0] matmult_out_b201,
    output wire signed [63:0] matmult_out_b202,
    output wire signed [63:0] matmult_out_b203,
    output wire signed [63:0] matmult_out_b204,
    output wire signed [63:0] matmult_out_b205,
    output wire signed [63:0] matmult_out_b206,
    output wire signed [63:0] matmult_out_b207,
    output wire signed [63:0] matmult_out_b208,
    output wire signed [63:0] matmult_out_b209,
    output wire signed [63:0] matmult_out_b210,
    output wire signed [63:0] matmult_out_b211,
    output wire signed [63:0] matmult_out_b212,
    output wire signed [63:0] matmult_out_b213,
    output wire signed [63:0] matmult_out_b214,
    output wire signed [63:0] matmult_out_b215,
    output wire signed [63:0] matmult_out_b216,
    output wire signed [63:0] matmult_out_b217,
    output wire signed [63:0] matmult_out_b218,
    output wire signed [63:0] matmult_out_b219,
    output wire signed [63:0] matmult_out_b220,
    output wire signed [63:0] matmult_out_b221,
    output wire signed [63:0] matmult_out_b222,
    output wire signed [63:0] matmult_out_b223,
    output wire signed [63:0] matmult_out_b224,
    output wire signed [63:0] matmult_out_b225,
    output wire signed [63:0] matmult_out_b226,
    output wire signed [63:0] matmult_out_b227,
    output wire signed [63:0] matmult_out_b228,
    output wire signed [63:0] matmult_out_b229,
    output wire signed [63:0] matmult_out_b230,
    output wire signed [63:0] matmult_out_b231,
    output wire signed [63:0] matmult_out_b232,
    output wire signed [63:0] matmult_out_b233,
    output wire signed [63:0] matmult_out_b234,
    output wire signed [63:0] matmult_out_b235,
    output wire signed [63:0] matmult_out_b236,
    output wire signed [63:0] matmult_out_b237,
    output wire signed [63:0] matmult_out_b238,
    output wire signed [63:0] matmult_out_b239,
    output wire signed [63:0] matmult_out_b240,
    output wire signed [63:0] matmult_out_b241,
    output wire signed [63:0] matmult_out_b242,
    output wire signed [63:0] matmult_out_b243,
    output wire signed [63:0] matmult_out_b244,
    output wire signed [63:0] matmult_out_b245,
    output wire signed [63:0] matmult_out_b246,
    output wire signed [63:0] matmult_out_b247,
    output wire signed [63:0] matmult_out_b248,
    output wire signed [63:0] matmult_out_b249,
    output wire signed [63:0] matmult_out_b250,
    output wire signed [63:0] matmult_out_b251,
    output wire signed [63:0] matmult_out_b252,
    output wire signed [63:0] matmult_out_b253,
    output wire signed [63:0] matmult_out_b254,
    output wire signed [63:0] matmult_out_b255,
    output wire signed [63:0] matmult_out_b256,
    output wire signed [63:0] matmult_out_b257,
    output wire signed [63:0] matmult_out_b258,
    output wire signed [63:0] matmult_out_b259,
    output wire signed [63:0] matmult_out_b260,
    output wire signed [63:0] matmult_out_b261,
    output wire signed [63:0] matmult_out_b262,
    output wire signed [63:0] matmult_out_b263,
    output wire signed [63:0] matmult_out_b264,
    output wire signed [63:0] matmult_out_b265,
    output wire signed [63:0] matmult_out_b266,
    output wire signed [63:0] matmult_out_b267,
    output wire signed [63:0] matmult_out_b268,
    output wire signed [63:0] matmult_out_b269,
    output wire signed [63:0] matmult_out_b270,
    output wire signed [63:0] matmult_out_b271,
    output wire signed [63:0] matmult_out_b272,
    output wire signed [63:0] matmult_out_b273,
    output wire signed [63:0] matmult_out_b274,
    output wire signed [63:0] matmult_out_b275,
    output wire signed [63:0] matmult_out_b276,
    output wire signed [63:0] matmult_out_b277,
    output wire signed [63:0] matmult_out_b278,
    output wire signed [63:0] matmult_out_b279,
    input wire [7:0] matmult_in_col,
    input wire signed [63:0] matmult_in_c0,
    input wire signed [63:0] matmult_in_c1,
    input wire signed [63:0] matmult_in_c2,
    input wire signed [63:0] matmult_in_c3,
    input wire signed [63:0] matmult_in_c4,
    input wire signed [63:0] matmult_in_c5,
    input wire signed [63:0] matmult_in_c6,
    input wire signed [63:0] matmult_in_c7,
    input wire signed [63:0] matmult_in_c8,
    input wire signed [63:0] matmult_in_c9,
    input wire signed [63:0] matmult_in_c10,
    input wire signed [63:0] matmult_in_c11,
    input wire signed [63:0] matmult_in_c12,
    input wire signed [63:0] matmult_in_c13,
    input wire signed [63:0] matmult_in_c14,
    input wire signed [63:0] matmult_in_c15,
    input wire signed [63:0] matmult_in_c16,
    input wire signed [63:0] matmult_in_c17,
    input wire signed [63:0] matmult_in_c18,
    input wire signed [63:0] matmult_in_c19,
    input wire signed [63:0] matmult_in_c20,
    input wire signed [63:0] matmult_in_c21,
    input wire signed [63:0] matmult_in_c22,
    input wire signed [63:0] matmult_in_c23,
    input wire signed [63:0] matmult_in_c24,
    input wire signed [63:0] matmult_in_c25,
    input wire signed [63:0] matmult_in_c26,
    input wire signed [63:0] matmult_in_c27,
    input wire signed [63:0] matmult_in_c28,
    input wire signed [63:0] matmult_in_c29,
    input wire signed [63:0] matmult_in_c30,
    input wire signed [63:0] matmult_in_c31,
    input wire signed [63:0] matmult_in_c32,
    input wire signed [63:0] matmult_in_c33,
    input wire signed [63:0] matmult_in_c34,
    input wire signed [63:0] matmult_in_c35,
    input wire signed [63:0] matmult_in_c36,
    input wire signed [63:0] matmult_in_c37,
    input wire signed [63:0] matmult_in_c38,
    input wire signed [63:0] matmult_in_c39,
    input wire signed [63:0] matmult_in_c40,
    input wire signed [63:0] matmult_in_c41,
    input wire signed [63:0] matmult_in_c42,
    input wire signed [63:0] matmult_in_c43,
    input wire signed [63:0] matmult_in_c44,
    input wire signed [63:0] matmult_in_c45,
    input wire signed [63:0] matmult_in_c46,
    input wire signed [63:0] matmult_in_c47,
    input wire signed [63:0] matmult_in_c48,
    input wire signed [63:0] matmult_in_c49,
    input wire signed [63:0] matmult_in_c50,
    input wire signed [63:0] matmult_in_c51,
    input wire signed [63:0] matmult_in_c52,
    input wire signed [63:0] matmult_in_c53,
    input wire signed [63:0] matmult_in_c54,
    input wire signed [63:0] matmult_in_c55,
    input wire signed [63:0] matmult_in_c56,
    input wire signed [63:0] matmult_in_c57,
    input wire signed [63:0] matmult_in_c58,
    input wire signed [63:0] matmult_in_c59,
    input wire signed [63:0] matmult_in_c60,
    input wire signed [63:0] matmult_in_c61,
    input wire signed [63:0] matmult_in_c62,
    input wire signed [63:0] matmult_in_c63,
    input wire signed [63:0] matmult_in_c64,
    input wire signed [63:0] matmult_in_c65,
    input wire signed [63:0] matmult_in_c66,
    input wire signed [63:0] matmult_in_c67,
    input wire signed [63:0] matmult_in_c68,
    input wire signed [63:0] matmult_in_c69,
    input wire signed [63:0] matmult_in_c70,
    input wire signed [63:0] matmult_in_c71,
    input wire signed [63:0] matmult_in_c72,
    input wire signed [63:0] matmult_in_c73,
    input wire signed [63:0] matmult_in_c74,
    input wire signed [63:0] matmult_in_c75,
    input wire signed [63:0] matmult_in_c76,
    input wire signed [63:0] matmult_in_c77,
    input wire signed [63:0] matmult_in_c78,
    input wire signed [63:0] matmult_in_c79,
    input wire signed [63:0] matmult_in_c80,
    input wire signed [63:0] matmult_in_c81,
    input wire signed [63:0] matmult_in_c82,
    input wire signed [63:0] matmult_in_c83,
    input wire signed [63:0] matmult_in_c84,
    input wire signed [63:0] matmult_in_c85,
    input wire signed [63:0] matmult_in_c86,
    input wire signed [63:0] matmult_in_c87,
    input wire signed [63:0] matmult_in_c88,
    input wire signed [63:0] matmult_in_c89,
    input wire signed [63:0] matmult_in_c90,
    input wire signed [63:0] matmult_in_c91,
    input wire signed [63:0] matmult_in_c92,
    input wire signed [63:0] matmult_in_c93,
    input wire signed [63:0] matmult_in_c94,
    input wire signed [63:0] matmult_in_c95,
    input wire signed [63:0] matmult_in_c96,
    input wire signed [63:0] matmult_in_c97,
    input wire signed [63:0] matmult_in_c98,
    input wire signed [63:0] matmult_in_c99,
    input wire signed [63:0] matmult_in_c100,
    input wire signed [63:0] matmult_in_c101,
    input wire signed [63:0] matmult_in_c102,
    input wire signed [63:0] matmult_in_c103,
    input wire signed [63:0] matmult_in_c104,
    input wire signed [63:0] matmult_in_c105,
    input wire signed [63:0] matmult_in_c106,
    input wire signed [63:0] matmult_in_c107,
    input wire signed [63:0] matmult_in_c108,
    input wire signed [63:0] matmult_in_c109,
    input wire signed [63:0] matmult_in_c110,
    input wire signed [63:0] matmult_in_c111,
    input wire signed [63:0] matmult_in_c112,
    input wire signed [63:0] matmult_in_c113,
    input wire signed [63:0] matmult_in_c114,
    input wire signed [63:0] matmult_in_c115,
    input wire signed [63:0] matmult_in_c116,
    input wire signed [63:0] matmult_in_c117,
    input wire signed [63:0] matmult_in_c118,
    input wire signed [63:0] matmult_in_c119,
    input wire signed [63:0] matmult_in_c120,
    input wire signed [63:0] matmult_in_c121,
    input wire signed [63:0] matmult_in_c122,
    input wire signed [63:0] matmult_in_c123,
    input wire signed [63:0] matmult_in_c124,
    input wire signed [63:0] matmult_in_c125,
    input wire signed [63:0] matmult_in_c126,
    input wire signed [63:0] matmult_in_c127,
    input wire signed [63:0] matmult_in_c128,
    input wire signed [63:0] matmult_in_c129,
    input wire signed [63:0] matmult_in_c130,
    input wire signed [63:0] matmult_in_c131,
    input wire signed [63:0] matmult_in_c132,
    input wire signed [63:0] matmult_in_c133,
    input wire signed [63:0] matmult_in_c134,
    input wire signed [63:0] matmult_in_c135,
    input wire signed [63:0] matmult_in_c136,
    input wire signed [63:0] matmult_in_c137,
    input wire signed [63:0] matmult_in_c138,
    input wire signed [63:0] matmult_in_c139,
    input wire signed [63:0] matmult_in_c140,
    input wire signed [63:0] matmult_in_c141,
    input wire signed [63:0] matmult_in_c142,
    input wire signed [63:0] matmult_in_c143,
    input wire signed [63:0] matmult_in_c144,
    input wire signed [63:0] matmult_in_c145,
    input wire signed [63:0] matmult_in_c146,
    input wire signed [63:0] matmult_in_c147,
    input wire signed [63:0] matmult_in_c148,
    input wire signed [63:0] matmult_in_c149,
    input wire signed [63:0] matmult_in_c150,
    input wire signed [63:0] matmult_in_c151,
    input wire signed [63:0] matmult_in_c152,
    input wire signed [63:0] matmult_in_c153,
    input wire signed [63:0] matmult_in_c154,
    input wire signed [63:0] matmult_in_c155,
    input wire signed [63:0] matmult_in_c156,
    input wire signed [63:0] matmult_in_c157,
    input wire signed [63:0] matmult_in_c158,
    input wire signed [63:0] matmult_in_c159,
    input wire signed [63:0] matmult_in_c160,
    input wire signed [63:0] matmult_in_c161,
    input wire signed [63:0] matmult_in_c162,
    input wire signed [63:0] matmult_in_c163,
    input wire signed [63:0] matmult_in_c164,
    input wire signed [63:0] matmult_in_c165,
    input wire signed [63:0] matmult_in_c166,
    input wire signed [63:0] matmult_in_c167,
    input wire signed [63:0] matmult_in_c168,
    input wire signed [63:0] matmult_in_c169,
    input wire signed [63:0] matmult_in_c170,
    input wire signed [63:0] matmult_in_c171,
    input wire signed [63:0] matmult_in_c172,
    input wire signed [63:0] matmult_in_c173,
    input wire signed [63:0] matmult_in_c174,
    input wire signed [63:0] matmult_in_c175,
    input wire signed [63:0] matmult_in_c176,
    input wire signed [63:0] matmult_in_c177,
    input wire signed [63:0] matmult_in_c178,
    input wire signed [63:0] matmult_in_c179,
    input wire signed [63:0] matmult_in_c180,
    input wire signed [63:0] matmult_in_c181,
    input wire signed [63:0] matmult_in_c182,
    input wire signed [63:0] matmult_in_c183,
    input wire signed [63:0] matmult_in_c184,
    input wire signed [63:0] matmult_in_c185,
    input wire signed [63:0] matmult_in_c186,
    input wire signed [63:0] matmult_in_c187,
    input wire signed [63:0] matmult_in_c188,
    input wire signed [63:0] matmult_in_c189,
    input wire signed [63:0] matmult_in_c190,
    input wire signed [63:0] matmult_in_c191,
    input wire signed [63:0] matmult_in_c192,
    input wire signed [63:0] matmult_in_c193,
    input wire signed [63:0] matmult_in_c194,
    input wire signed [63:0] matmult_in_c195,
    input wire signed [63:0] matmult_in_c196,
    input wire signed [63:0] matmult_in_c197,
    input wire signed [63:0] matmult_in_c198,
    input wire signed [63:0] matmult_in_c199,
    input wire signed [63:0] matmult_in_c200,
    input wire signed [63:0] matmult_in_c201,
    input wire signed [63:0] matmult_in_c202,
    input wire signed [63:0] matmult_in_c203,
    input wire signed [63:0] matmult_in_c204,
    input wire signed [63:0] matmult_in_c205,
    input wire signed [63:0] matmult_in_c206,
    input wire signed [63:0] matmult_in_c207,
    input wire signed [63:0] matmult_in_c208,
    input wire signed [63:0] matmult_in_c209,
    input wire signed [63:0] matmult_in_c210,
    input wire signed [63:0] matmult_in_c211,
    input wire signed [63:0] matmult_in_c212,
    input wire signed [63:0] matmult_in_c213,
    input wire signed [63:0] matmult_in_c214,
    input wire signed [63:0] matmult_in_c215,
    input wire signed [63:0] matmult_in_c216,
    input wire signed [63:0] matmult_in_c217,
    input wire signed [63:0] matmult_in_c218,
    input wire signed [63:0] matmult_in_c219,
    input wire signed [63:0] matmult_in_c220,
    input wire signed [63:0] matmult_in_c221,
    input wire signed [63:0] matmult_in_c222,
    input wire signed [63:0] matmult_in_c223,
    input wire signed [63:0] matmult_in_c224,
    input wire signed [63:0] matmult_in_c225,
    input wire signed [63:0] matmult_in_c226,
    input wire signed [63:0] matmult_in_c227,
    input wire signed [63:0] matmult_in_c228,
    input wire signed [63:0] matmult_in_c229,
    input wire signed [63:0] matmult_in_c230,
    input wire signed [63:0] matmult_in_c231,
    input wire signed [63:0] matmult_in_c232,
    input wire signed [63:0] matmult_in_c233,
    input wire signed [63:0] matmult_in_c234,
    input wire signed [63:0] matmult_in_c235,
    input wire signed [63:0] matmult_in_c236,
    input wire signed [63:0] matmult_in_c237,
    input wire signed [63:0] matmult_in_c238,
    input wire signed [63:0] matmult_in_c239,
    input wire signed [63:0] matmult_in_c240,
    input wire signed [63:0] matmult_in_c241,
    input wire signed [63:0] matmult_in_c242,
    input wire signed [63:0] matmult_in_c243,
    input wire signed [63:0] matmult_in_c244,
    input wire signed [63:0] matmult_in_c245,
    input wire signed [63:0] matmult_in_c246,
    input wire signed [63:0] matmult_in_c247,
    input wire signed [63:0] matmult_in_c248,
    input wire signed [63:0] matmult_in_c249,
    input wire signed [63:0] matmult_in_c250,
    input wire signed [63:0] matmult_in_c251,
    input wire signed [63:0] matmult_in_c252,
    input wire signed [63:0] matmult_in_c253,
    input wire signed [63:0] matmult_in_c254,
    input wire signed [63:0] matmult_in_c255,
    input wire signed [63:0] matmult_in_c256,
    input wire signed [63:0] matmult_in_c257,
    input wire signed [63:0] matmult_in_c258,
    input wire signed [63:0] matmult_in_c259,
    input wire signed [63:0] matmult_in_c260,
    input wire signed [63:0] matmult_in_c261,
    input wire signed [63:0] matmult_in_c262,
    input wire signed [63:0] matmult_in_c263,
    input wire signed [63:0] matmult_in_c264,
    input wire signed [63:0] matmult_in_c265,
    input wire signed [63:0] matmult_in_c266,
    input wire signed [63:0] matmult_in_c267,
    input wire signed [63:0] matmult_in_c268,
    input wire signed [63:0] matmult_in_c269,
    input wire signed [63:0] matmult_in_c270,
    input wire signed [63:0] matmult_in_c271,
    input wire signed [63:0] matmult_in_c272,
    input wire signed [63:0] matmult_in_c273,
    input wire signed [63:0] matmult_in_c274,
    input wire signed [63:0] matmult_in_c275,
    input wire signed [63:0] matmult_in_c276,
    input wire signed [63:0] matmult_in_c277,
    input wire signed [63:0] matmult_in_c278,
    input wire signed [63:0] matmult_in_c279,
    output wire signed [63:0] matmult_out_c0,
    output wire signed [63:0] matmult_out_c1,
    output wire signed [63:0] matmult_out_c2,
    output wire signed [63:0] matmult_out_c3,
    output wire signed [63:0] matmult_out_c4,
    output wire signed [63:0] matmult_out_c5,
    output wire signed [63:0] matmult_out_c6,
    output wire signed [63:0] matmult_out_c7,
    output wire signed [63:0] matmult_out_c8,
    output wire signed [63:0] matmult_out_c9,
    output wire signed [63:0] matmult_out_c10,
    output wire signed [63:0] matmult_out_c11,
    output wire signed [63:0] matmult_out_c12,
    output wire signed [63:0] matmult_out_c13,
    output wire signed [63:0] matmult_out_c14,
    output wire signed [63:0] matmult_out_c15,
    output wire signed [63:0] matmult_out_c16,
    output wire signed [63:0] matmult_out_c17,
    output wire signed [63:0] matmult_out_c18,
    output wire signed [63:0] matmult_out_c19,
    output wire signed [63:0] matmult_out_c20,
    output wire signed [63:0] matmult_out_c21,
    output wire signed [63:0] matmult_out_c22,
    output wire signed [63:0] matmult_out_c23,
    output wire signed [63:0] matmult_out_c24,
    output wire signed [63:0] matmult_out_c25,
    output wire signed [63:0] matmult_out_c26,
    output wire signed [63:0] matmult_out_c27,
    output wire signed [63:0] matmult_out_c28,
    output wire signed [63:0] matmult_out_c29,
    output wire signed [63:0] matmult_out_c30,
    output wire signed [63:0] matmult_out_c31,
    output wire signed [63:0] matmult_out_c32,
    output wire signed [63:0] matmult_out_c33,
    output wire signed [63:0] matmult_out_c34,
    output wire signed [63:0] matmult_out_c35,
    output wire signed [63:0] matmult_out_c36,
    output wire signed [63:0] matmult_out_c37,
    output wire signed [63:0] matmult_out_c38,
    output wire signed [63:0] matmult_out_c39,
    output wire signed [63:0] matmult_out_c40,
    output wire signed [63:0] matmult_out_c41,
    output wire signed [63:0] matmult_out_c42,
    output wire signed [63:0] matmult_out_c43,
    output wire signed [63:0] matmult_out_c44,
    output wire signed [63:0] matmult_out_c45,
    output wire signed [63:0] matmult_out_c46,
    output wire signed [63:0] matmult_out_c47,
    output wire signed [63:0] matmult_out_c48,
    output wire signed [63:0] matmult_out_c49,
    output wire signed [63:0] matmult_out_c50,
    output wire signed [63:0] matmult_out_c51,
    output wire signed [63:0] matmult_out_c52,
    output wire signed [63:0] matmult_out_c53,
    output wire signed [63:0] matmult_out_c54,
    output wire signed [63:0] matmult_out_c55,
    output wire signed [63:0] matmult_out_c56,
    output wire signed [63:0] matmult_out_c57,
    output wire signed [63:0] matmult_out_c58,
    output wire signed [63:0] matmult_out_c59,
    output wire signed [63:0] matmult_out_c60,
    output wire signed [63:0] matmult_out_c61,
    output wire signed [63:0] matmult_out_c62,
    output wire signed [63:0] matmult_out_c63,
    output wire signed [63:0] matmult_out_c64,
    output wire signed [63:0] matmult_out_c65,
    output wire signed [63:0] matmult_out_c66,
    output wire signed [63:0] matmult_out_c67,
    output wire signed [63:0] matmult_out_c68,
    output wire signed [63:0] matmult_out_c69,
    output wire signed [63:0] matmult_out_c70,
    output wire signed [63:0] matmult_out_c71,
    output wire signed [63:0] matmult_out_c72,
    output wire signed [63:0] matmult_out_c73,
    output wire signed [63:0] matmult_out_c74,
    output wire signed [63:0] matmult_out_c75,
    output wire signed [63:0] matmult_out_c76,
    output wire signed [63:0] matmult_out_c77,
    output wire signed [63:0] matmult_out_c78,
    output wire signed [63:0] matmult_out_c79,
    output wire signed [63:0] matmult_out_c80,
    output wire signed [63:0] matmult_out_c81,
    output wire signed [63:0] matmult_out_c82,
    output wire signed [63:0] matmult_out_c83,
    output wire signed [63:0] matmult_out_c84,
    output wire signed [63:0] matmult_out_c85,
    output wire signed [63:0] matmult_out_c86,
    output wire signed [63:0] matmult_out_c87,
    output wire signed [63:0] matmult_out_c88,
    output wire signed [63:0] matmult_out_c89,
    output wire signed [63:0] matmult_out_c90,
    output wire signed [63:0] matmult_out_c91,
    output wire signed [63:0] matmult_out_c92,
    output wire signed [63:0] matmult_out_c93,
    output wire signed [63:0] matmult_out_c94,
    output wire signed [63:0] matmult_out_c95,
    output wire signed [63:0] matmult_out_c96,
    output wire signed [63:0] matmult_out_c97,
    output wire signed [63:0] matmult_out_c98,
    output wire signed [63:0] matmult_out_c99,
    output wire signed [63:0] matmult_out_c100,
    output wire signed [63:0] matmult_out_c101,
    output wire signed [63:0] matmult_out_c102,
    output wire signed [63:0] matmult_out_c103,
    output wire signed [63:0] matmult_out_c104,
    output wire signed [63:0] matmult_out_c105,
    output wire signed [63:0] matmult_out_c106,
    output wire signed [63:0] matmult_out_c107,
    output wire signed [63:0] matmult_out_c108,
    output wire signed [63:0] matmult_out_c109,
    output wire signed [63:0] matmult_out_c110,
    output wire signed [63:0] matmult_out_c111,
    output wire signed [63:0] matmult_out_c112,
    output wire signed [63:0] matmult_out_c113,
    output wire signed [63:0] matmult_out_c114,
    output wire signed [63:0] matmult_out_c115,
    output wire signed [63:0] matmult_out_c116,
    output wire signed [63:0] matmult_out_c117,
    output wire signed [63:0] matmult_out_c118,
    output wire signed [63:0] matmult_out_c119,
    output wire signed [63:0] matmult_out_c120,
    output wire signed [63:0] matmult_out_c121,
    output wire signed [63:0] matmult_out_c122,
    output wire signed [63:0] matmult_out_c123,
    output wire signed [63:0] matmult_out_c124,
    output wire signed [63:0] matmult_out_c125,
    output wire signed [63:0] matmult_out_c126,
    output wire signed [63:0] matmult_out_c127,
    output wire signed [63:0] matmult_out_c128,
    output wire signed [63:0] matmult_out_c129,
    output wire signed [63:0] matmult_out_c130,
    output wire signed [63:0] matmult_out_c131,
    output wire signed [63:0] matmult_out_c132,
    output wire signed [63:0] matmult_out_c133,
    output wire signed [63:0] matmult_out_c134,
    output wire signed [63:0] matmult_out_c135,
    output wire signed [63:0] matmult_out_c136,
    output wire signed [63:0] matmult_out_c137,
    output wire signed [63:0] matmult_out_c138,
    output wire signed [63:0] matmult_out_c139,
    output wire signed [63:0] matmult_out_c140,
    output wire signed [63:0] matmult_out_c141,
    output wire signed [63:0] matmult_out_c142,
    output wire signed [63:0] matmult_out_c143,
    output wire signed [63:0] matmult_out_c144,
    output wire signed [63:0] matmult_out_c145,
    output wire signed [63:0] matmult_out_c146,
    output wire signed [63:0] matmult_out_c147,
    output wire signed [63:0] matmult_out_c148,
    output wire signed [63:0] matmult_out_c149,
    output wire signed [63:0] matmult_out_c150,
    output wire signed [63:0] matmult_out_c151,
    output wire signed [63:0] matmult_out_c152,
    output wire signed [63:0] matmult_out_c153,
    output wire signed [63:0] matmult_out_c154,
    output wire signed [63:0] matmult_out_c155,
    output wire signed [63:0] matmult_out_c156,
    output wire signed [63:0] matmult_out_c157,
    output wire signed [63:0] matmult_out_c158,
    output wire signed [63:0] matmult_out_c159,
    output wire signed [63:0] matmult_out_c160,
    output wire signed [63:0] matmult_out_c161,
    output wire signed [63:0] matmult_out_c162,
    output wire signed [63:0] matmult_out_c163,
    output wire signed [63:0] matmult_out_c164,
    output wire signed [63:0] matmult_out_c165,
    output wire signed [63:0] matmult_out_c166,
    output wire signed [63:0] matmult_out_c167,
    output wire signed [63:0] matmult_out_c168,
    output wire signed [63:0] matmult_out_c169,
    output wire signed [63:0] matmult_out_c170,
    output wire signed [63:0] matmult_out_c171,
    output wire signed [63:0] matmult_out_c172,
    output wire signed [63:0] matmult_out_c173,
    output wire signed [63:0] matmult_out_c174,
    output wire signed [63:0] matmult_out_c175,
    output wire signed [63:0] matmult_out_c176,
    output wire signed [63:0] matmult_out_c177,
    output wire signed [63:0] matmult_out_c178,
    output wire signed [63:0] matmult_out_c179,
    output wire signed [63:0] matmult_out_c180,
    output wire signed [63:0] matmult_out_c181,
    output wire signed [63:0] matmult_out_c182,
    output wire signed [63:0] matmult_out_c183,
    output wire signed [63:0] matmult_out_c184,
    output wire signed [63:0] matmult_out_c185,
    output wire signed [63:0] matmult_out_c186,
    output wire signed [63:0] matmult_out_c187,
    output wire signed [63:0] matmult_out_c188,
    output wire signed [63:0] matmult_out_c189,
    output wire signed [63:0] matmult_out_c190,
    output wire signed [63:0] matmult_out_c191,
    output wire signed [63:0] matmult_out_c192,
    output wire signed [63:0] matmult_out_c193,
    output wire signed [63:0] matmult_out_c194,
    output wire signed [63:0] matmult_out_c195,
    output wire signed [63:0] matmult_out_c196,
    output wire signed [63:0] matmult_out_c197,
    output wire signed [63:0] matmult_out_c198,
    output wire signed [63:0] matmult_out_c199,
    output wire signed [63:0] matmult_out_c200,
    output wire signed [63:0] matmult_out_c201,
    output wire signed [63:0] matmult_out_c202,
    output wire signed [63:0] matmult_out_c203,
    output wire signed [63:0] matmult_out_c204,
    output wire signed [63:0] matmult_out_c205,
    output wire signed [63:0] matmult_out_c206,
    output wire signed [63:0] matmult_out_c207,
    output wire signed [63:0] matmult_out_c208,
    output wire signed [63:0] matmult_out_c209,
    output wire signed [63:0] matmult_out_c210,
    output wire signed [63:0] matmult_out_c211,
    output wire signed [63:0] matmult_out_c212,
    output wire signed [63:0] matmult_out_c213,
    output wire signed [63:0] matmult_out_c214,
    output wire signed [63:0] matmult_out_c215,
    output wire signed [63:0] matmult_out_c216,
    output wire signed [63:0] matmult_out_c217,
    output wire signed [63:0] matmult_out_c218,
    output wire signed [63:0] matmult_out_c219,
    output wire signed [63:0] matmult_out_c220,
    output wire signed [63:0] matmult_out_c221,
    output wire signed [63:0] matmult_out_c222,
    output wire signed [63:0] matmult_out_c223,
    output wire signed [63:0] matmult_out_c224,
    output wire signed [63:0] matmult_out_c225,
    output wire signed [63:0] matmult_out_c226,
    output wire signed [63:0] matmult_out_c227,
    output wire signed [63:0] matmult_out_c228,
    output wire signed [63:0] matmult_out_c229,
    output wire signed [63:0] matmult_out_c230,
    output wire signed [63:0] matmult_out_c231,
    output wire signed [63:0] matmult_out_c232,
    output wire signed [63:0] matmult_out_c233,
    output wire signed [63:0] matmult_out_c234,
    output wire signed [63:0] matmult_out_c235,
    output wire signed [63:0] matmult_out_c236,
    output wire signed [63:0] matmult_out_c237,
    output wire signed [63:0] matmult_out_c238,
    output wire signed [63:0] matmult_out_c239,
    output wire signed [63:0] matmult_out_c240,
    output wire signed [63:0] matmult_out_c241,
    output wire signed [63:0] matmult_out_c242,
    output wire signed [63:0] matmult_out_c243,
    output wire signed [63:0] matmult_out_c244,
    output wire signed [63:0] matmult_out_c245,
    output wire signed [63:0] matmult_out_c246,
    output wire signed [63:0] matmult_out_c247,
    output wire signed [63:0] matmult_out_c248,
    output wire signed [63:0] matmult_out_c249,
    output wire signed [63:0] matmult_out_c250,
    output wire signed [63:0] matmult_out_c251,
    output wire signed [63:0] matmult_out_c252,
    output wire signed [63:0] matmult_out_c253,
    output wire signed [63:0] matmult_out_c254,
    output wire signed [63:0] matmult_out_c255,
    output wire signed [63:0] matmult_out_c256,
    output wire signed [63:0] matmult_out_c257,
    output wire signed [63:0] matmult_out_c258,
    output wire signed [63:0] matmult_out_c259,
    output wire signed [63:0] matmult_out_c260,
    output wire signed [63:0] matmult_out_c261,
    output wire signed [63:0] matmult_out_c262,
    output wire signed [63:0] matmult_out_c263,
    output wire signed [63:0] matmult_out_c264,
    output wire signed [63:0] matmult_out_c265,
    output wire signed [63:0] matmult_out_c266,
    output wire signed [63:0] matmult_out_c267,
    output wire signed [63:0] matmult_out_c268,
    output wire signed [63:0] matmult_out_c269,
    output wire signed [63:0] matmult_out_c270,
    output wire signed [63:0] matmult_out_c271,
    output wire signed [63:0] matmult_out_c272,
    output wire signed [63:0] matmult_out_c273,
    output wire signed [63:0] matmult_out_c274,
    output wire signed [63:0] matmult_out_c275,
    output wire signed [63:0] matmult_out_c276,
    output wire signed [63:0] matmult_out_c277,
    output wire signed [63:0] matmult_out_c278,
    output wire signed [63:0] matmult_out_c279
);
    localparam idle = 0;
    localparam fin = 1;
    localparam calc = 2;
    reg [63:0] a[0:279];
    reg [63:0] b[0:279];
    reg [63:0] c[0:279];
    reg [1:0] state;

    assign matmult_out_c0 = c[0];
    assign matmult_out_c1 = c[1];
    assign matmult_out_c2 = c[2];
    assign matmult_out_c3 = c[3];
    assign matmult_out_c4 = c[4];
    assign matmult_out_c5 = c[5];
    assign matmult_out_c6 = c[6];
    assign matmult_out_c7 = c[7];
    assign matmult_out_c8 = c[8];
    assign matmult_out_c9 = c[9];
    assign matmult_out_c10 = c[10];
    assign matmult_out_c11 = c[11];
    assign matmult_out_c12 = c[12];
    assign matmult_out_c13 = c[13];
    assign matmult_out_c14 = c[14];
    assign matmult_out_c15 = c[15];
    assign matmult_out_c16 = c[16];
    assign matmult_out_c17 = c[17];
    assign matmult_out_c18 = c[18];
    assign matmult_out_c19 = c[19];
    assign matmult_out_c20 = c[20];
    assign matmult_out_c21 = c[21];
    assign matmult_out_c22 = c[22];
    assign matmult_out_c23 = c[23];
    assign matmult_out_c24 = c[24];
    assign matmult_out_c25 = c[25];
    assign matmult_out_c26 = c[26];
    assign matmult_out_c27 = c[27];
    assign matmult_out_c28 = c[28];
    assign matmult_out_c29 = c[29];
    assign matmult_out_c30 = c[30];
    assign matmult_out_c31 = c[31];
    assign matmult_out_c32 = c[32];
    assign matmult_out_c33 = c[33];
    assign matmult_out_c34 = c[34];
    assign matmult_out_c35 = c[35];
    assign matmult_out_c36 = c[36];
    assign matmult_out_c37 = c[37];
    assign matmult_out_c38 = c[38];
    assign matmult_out_c39 = c[39];
    assign matmult_out_c40 = c[40];
    assign matmult_out_c41 = c[41];
    assign matmult_out_c42 = c[42];
    assign matmult_out_c43 = c[43];
    assign matmult_out_c44 = c[44];
    assign matmult_out_c45 = c[45];
    assign matmult_out_c46 = c[46];
    assign matmult_out_c47 = c[47];
    assign matmult_out_c48 = c[48];
    assign matmult_out_c49 = c[49];
    assign matmult_out_c50 = c[50];
    assign matmult_out_c51 = c[51];
    assign matmult_out_c52 = c[52];
    assign matmult_out_c53 = c[53];
    assign matmult_out_c54 = c[54];
    assign matmult_out_c55 = c[55];
    assign matmult_out_c56 = c[56];
    assign matmult_out_c57 = c[57];
    assign matmult_out_c58 = c[58];
    assign matmult_out_c59 = c[59];
    assign matmult_out_c60 = c[60];
    assign matmult_out_c61 = c[61];
    assign matmult_out_c62 = c[62];
    assign matmult_out_c63 = c[63];
    assign matmult_out_c64 = c[64];
    assign matmult_out_c65 = c[65];
    assign matmult_out_c66 = c[66];
    assign matmult_out_c67 = c[67];
    assign matmult_out_c68 = c[68];
    assign matmult_out_c69 = c[69];
    assign matmult_out_c70 = c[70];
    assign matmult_out_c71 = c[71];
    assign matmult_out_c72 = c[72];
    assign matmult_out_c73 = c[73];
    assign matmult_out_c74 = c[74];
    assign matmult_out_c75 = c[75];
    assign matmult_out_c76 = c[76];
    assign matmult_out_c77 = c[77];
    assign matmult_out_c78 = c[78];
    assign matmult_out_c79 = c[79];
    assign matmult_out_c80 = c[80];
    assign matmult_out_c81 = c[81];
    assign matmult_out_c82 = c[82];
    assign matmult_out_c83 = c[83];
    assign matmult_out_c84 = c[84];
    assign matmult_out_c85 = c[85];
    assign matmult_out_c86 = c[86];
    assign matmult_out_c87 = c[87];
    assign matmult_out_c88 = c[88];
    assign matmult_out_c89 = c[89];
    assign matmult_out_c90 = c[90];
    assign matmult_out_c91 = c[91];
    assign matmult_out_c92 = c[92];
    assign matmult_out_c93 = c[93];
    assign matmult_out_c94 = c[94];
    assign matmult_out_c95 = c[95];
    assign matmult_out_c96 = c[96];
    assign matmult_out_c97 = c[97];
    assign matmult_out_c98 = c[98];
    assign matmult_out_c99 = c[99];
    assign matmult_out_c100 = c[100];
    assign matmult_out_c101 = c[101];
    assign matmult_out_c102 = c[102];
    assign matmult_out_c103 = c[103];
    assign matmult_out_c104 = c[104];
    assign matmult_out_c105 = c[105];
    assign matmult_out_c106 = c[106];
    assign matmult_out_c107 = c[107];
    assign matmult_out_c108 = c[108];
    assign matmult_out_c109 = c[109];
    assign matmult_out_c110 = c[110];
    assign matmult_out_c111 = c[111];
    assign matmult_out_c112 = c[112];
    assign matmult_out_c113 = c[113];
    assign matmult_out_c114 = c[114];
    assign matmult_out_c115 = c[115];
    assign matmult_out_c116 = c[116];
    assign matmult_out_c117 = c[117];
    assign matmult_out_c118 = c[118];
    assign matmult_out_c119 = c[119];
    assign matmult_out_c120 = c[120];
    assign matmult_out_c121 = c[121];
    assign matmult_out_c122 = c[122];
    assign matmult_out_c123 = c[123];
    assign matmult_out_c124 = c[124];
    assign matmult_out_c125 = c[125];
    assign matmult_out_c126 = c[126];
    assign matmult_out_c127 = c[127];
    assign matmult_out_c128 = c[128];
    assign matmult_out_c129 = c[129];
    assign matmult_out_c130 = c[130];
    assign matmult_out_c131 = c[131];
    assign matmult_out_c132 = c[132];
    assign matmult_out_c133 = c[133];
    assign matmult_out_c134 = c[134];
    assign matmult_out_c135 = c[135];
    assign matmult_out_c136 = c[136];
    assign matmult_out_c137 = c[137];
    assign matmult_out_c138 = c[138];
    assign matmult_out_c139 = c[139];
    assign matmult_out_c140 = c[140];
    assign matmult_out_c141 = c[141];
    assign matmult_out_c142 = c[142];
    assign matmult_out_c143 = c[143];
    assign matmult_out_c144 = c[144];
    assign matmult_out_c145 = c[145];
    assign matmult_out_c146 = c[146];
    assign matmult_out_c147 = c[147];
    assign matmult_out_c148 = c[148];
    assign matmult_out_c149 = c[149];
    assign matmult_out_c150 = c[150];
    assign matmult_out_c151 = c[151];
    assign matmult_out_c152 = c[152];
    assign matmult_out_c153 = c[153];
    assign matmult_out_c154 = c[154];
    assign matmult_out_c155 = c[155];
    assign matmult_out_c156 = c[156];
    assign matmult_out_c157 = c[157];
    assign matmult_out_c158 = c[158];
    assign matmult_out_c159 = c[159];
    assign matmult_out_c160 = c[160];
    assign matmult_out_c161 = c[161];
    assign matmult_out_c162 = c[162];
    assign matmult_out_c163 = c[163];
    assign matmult_out_c164 = c[164];
    assign matmult_out_c165 = c[165];
    assign matmult_out_c166 = c[166];
    assign matmult_out_c167 = c[167];
    assign matmult_out_c168 = c[168];
    assign matmult_out_c169 = c[169];
    assign matmult_out_c170 = c[170];
    assign matmult_out_c171 = c[171];
    assign matmult_out_c172 = c[172];
    assign matmult_out_c173 = c[173];
    assign matmult_out_c174 = c[174];
    assign matmult_out_c175 = c[175];
    assign matmult_out_c176 = c[176];
    assign matmult_out_c177 = c[177];
    assign matmult_out_c178 = c[178];
    assign matmult_out_c179 = c[179];
    assign matmult_out_c180 = c[180];
    assign matmult_out_c181 = c[181];
    assign matmult_out_c182 = c[182];
    assign matmult_out_c183 = c[183];
    assign matmult_out_c184 = c[184];
    assign matmult_out_c185 = c[185];
    assign matmult_out_c186 = c[186];
    assign matmult_out_c187 = c[187];
    assign matmult_out_c188 = c[188];
    assign matmult_out_c189 = c[189];
    assign matmult_out_c190 = c[190];
    assign matmult_out_c191 = c[191];
    assign matmult_out_c192 = c[192];
    assign matmult_out_c193 = c[193];
    assign matmult_out_c194 = c[194];
    assign matmult_out_c195 = c[195];
    assign matmult_out_c196 = c[196];
    assign matmult_out_c197 = c[197];
    assign matmult_out_c198 = c[198];
    assign matmult_out_c199 = c[199];
    assign matmult_out_c200 = c[200];
    assign matmult_out_c201 = c[201];
    assign matmult_out_c202 = c[202];
    assign matmult_out_c203 = c[203];
    assign matmult_out_c204 = c[204];
    assign matmult_out_c205 = c[205];
    assign matmult_out_c206 = c[206];
    assign matmult_out_c207 = c[207];
    assign matmult_out_c208 = c[208];
    assign matmult_out_c209 = c[209];
    assign matmult_out_c210 = c[210];
    assign matmult_out_c211 = c[211];
    assign matmult_out_c212 = c[212];
    assign matmult_out_c213 = c[213];
    assign matmult_out_c214 = c[214];
    assign matmult_out_c215 = c[215];
    assign matmult_out_c216 = c[216];
    assign matmult_out_c217 = c[217];
    assign matmult_out_c218 = c[218];
    assign matmult_out_c219 = c[219];
    assign matmult_out_c220 = c[220];
    assign matmult_out_c221 = c[221];
    assign matmult_out_c222 = c[222];
    assign matmult_out_c223 = c[223];
    assign matmult_out_c224 = c[224];
    assign matmult_out_c225 = c[225];
    assign matmult_out_c226 = c[226];
    assign matmult_out_c227 = c[227];
    assign matmult_out_c228 = c[228];
    assign matmult_out_c229 = c[229];
    assign matmult_out_c230 = c[230];
    assign matmult_out_c231 = c[231];
    assign matmult_out_c232 = c[232];
    assign matmult_out_c233 = c[233];
    assign matmult_out_c234 = c[234];
    assign matmult_out_c235 = c[235];
    assign matmult_out_c236 = c[236];
    assign matmult_out_c237 = c[237];
    assign matmult_out_c238 = c[238];
    assign matmult_out_c239 = c[239];
    assign matmult_out_c240 = c[240];
    assign matmult_out_c241 = c[241];
    assign matmult_out_c242 = c[242];
    assign matmult_out_c243 = c[243];
    assign matmult_out_c244 = c[244];
    assign matmult_out_c245 = c[245];
    assign matmult_out_c246 = c[246];
    assign matmult_out_c247 = c[247];
    assign matmult_out_c248 = c[248];
    assign matmult_out_c249 = c[249];
    assign matmult_out_c250 = c[250];
    assign matmult_out_c251 = c[251];
    assign matmult_out_c252 = c[252];
    assign matmult_out_c253 = c[253];
    assign matmult_out_c254 = c[254];
    assign matmult_out_c255 = c[255];
    assign matmult_out_c256 = c[256];
    assign matmult_out_c257 = c[257];
    assign matmult_out_c258 = c[258];
    assign matmult_out_c259 = c[259];
    assign matmult_out_c260 = c[260];
    assign matmult_out_c261 = c[261];
    assign matmult_out_c262 = c[262];
    assign matmult_out_c263 = c[263];
    assign matmult_out_c264 = c[264];
    assign matmult_out_c265 = c[265];
    assign matmult_out_c266 = c[266];
    assign matmult_out_c267 = c[267];
    assign matmult_out_c268 = c[268];
    assign matmult_out_c269 = c[269];
    assign matmult_out_c270 = c[270];
    assign matmult_out_c271 = c[271];
    assign matmult_out_c272 = c[272];
    assign matmult_out_c273 = c[273];
    assign matmult_out_c274 = c[274];
    assign matmult_out_c275 = c[275];
    assign matmult_out_c276 = c[276];
    assign matmult_out_c277 = c[277];
    assign matmult_out_c278 = c[278];
    assign matmult_out_c279 = c[279];

    always @(posedge clk) begin
        if (rst) begin
            for (integer i = 0; i < 280; i++) begin
    a[i] <= 0;
end
            for (integer i = 0; i < 280; i++) begin
    b[i] <= 0;
end
            for (integer i = 0; i < 280; i++) begin
    c[i] <= 0;
end
            state <= 0;
            matmult_valid <= 0;
        end else begin
            case (state)
                idle: begin
                    matmult_valid <= 0;
                    if (matmult_ready) begin
    a[0] <= matmult_in_a0;
    a[1] <= matmult_in_a1;
    a[2] <= matmult_in_a2;
    a[3] <= matmult_in_a3;
    a[4] <= matmult_in_a4;
    a[5] <= matmult_in_a5;
    a[6] <= matmult_in_a6;
    a[7] <= matmult_in_a7;
    a[8] <= matmult_in_a8;
    a[9] <= matmult_in_a9;
    a[10] <= matmult_in_a10;
    a[11] <= matmult_in_a11;
    a[12] <= matmult_in_a12;
    a[13] <= matmult_in_a13;
    a[14] <= matmult_in_a14;
    a[15] <= matmult_in_a15;
    a[16] <= matmult_in_a16;
    a[17] <= matmult_in_a17;
    a[18] <= matmult_in_a18;
    a[19] <= matmult_in_a19;
    a[20] <= matmult_in_a20;
    a[21] <= matmult_in_a21;
    a[22] <= matmult_in_a22;
    a[23] <= matmult_in_a23;
    a[24] <= matmult_in_a24;
    a[25] <= matmult_in_a25;
    a[26] <= matmult_in_a26;
    a[27] <= matmult_in_a27;
    a[28] <= matmult_in_a28;
    a[29] <= matmult_in_a29;
    a[30] <= matmult_in_a30;
    a[31] <= matmult_in_a31;
    a[32] <= matmult_in_a32;
    a[33] <= matmult_in_a33;
    a[34] <= matmult_in_a34;
    a[35] <= matmult_in_a35;
    a[36] <= matmult_in_a36;
    a[37] <= matmult_in_a37;
    a[38] <= matmult_in_a38;
    a[39] <= matmult_in_a39;
    a[40] <= matmult_in_a40;
    a[41] <= matmult_in_a41;
    a[42] <= matmult_in_a42;
    a[43] <= matmult_in_a43;
    a[44] <= matmult_in_a44;
    a[45] <= matmult_in_a45;
    a[46] <= matmult_in_a46;
    a[47] <= matmult_in_a47;
    a[48] <= matmult_in_a48;
    a[49] <= matmult_in_a49;
    a[50] <= matmult_in_a50;
    a[51] <= matmult_in_a51;
    a[52] <= matmult_in_a52;
    a[53] <= matmult_in_a53;
    a[54] <= matmult_in_a54;
    a[55] <= matmult_in_a55;
    a[56] <= matmult_in_a56;
    a[57] <= matmult_in_a57;
    a[58] <= matmult_in_a58;
    a[59] <= matmult_in_a59;
    a[60] <= matmult_in_a60;
    a[61] <= matmult_in_a61;
    a[62] <= matmult_in_a62;
    a[63] <= matmult_in_a63;
    a[64] <= matmult_in_a64;
    a[65] <= matmult_in_a65;
    a[66] <= matmult_in_a66;
    a[67] <= matmult_in_a67;
    a[68] <= matmult_in_a68;
    a[69] <= matmult_in_a69;
    a[70] <= matmult_in_a70;
    a[71] <= matmult_in_a71;
    a[72] <= matmult_in_a72;
    a[73] <= matmult_in_a73;
    a[74] <= matmult_in_a74;
    a[75] <= matmult_in_a75;
    a[76] <= matmult_in_a76;
    a[77] <= matmult_in_a77;
    a[78] <= matmult_in_a78;
    a[79] <= matmult_in_a79;
    a[80] <= matmult_in_a80;
    a[81] <= matmult_in_a81;
    a[82] <= matmult_in_a82;
    a[83] <= matmult_in_a83;
    a[84] <= matmult_in_a84;
    a[85] <= matmult_in_a85;
    a[86] <= matmult_in_a86;
    a[87] <= matmult_in_a87;
    a[88] <= matmult_in_a88;
    a[89] <= matmult_in_a89;
    a[90] <= matmult_in_a90;
    a[91] <= matmult_in_a91;
    a[92] <= matmult_in_a92;
    a[93] <= matmult_in_a93;
    a[94] <= matmult_in_a94;
    a[95] <= matmult_in_a95;
    a[96] <= matmult_in_a96;
    a[97] <= matmult_in_a97;
    a[98] <= matmult_in_a98;
    a[99] <= matmult_in_a99;
    a[100] <= matmult_in_a100;
    a[101] <= matmult_in_a101;
    a[102] <= matmult_in_a102;
    a[103] <= matmult_in_a103;
    a[104] <= matmult_in_a104;
    a[105] <= matmult_in_a105;
    a[106] <= matmult_in_a106;
    a[107] <= matmult_in_a107;
    a[108] <= matmult_in_a108;
    a[109] <= matmult_in_a109;
    a[110] <= matmult_in_a110;
    a[111] <= matmult_in_a111;
    a[112] <= matmult_in_a112;
    a[113] <= matmult_in_a113;
    a[114] <= matmult_in_a114;
    a[115] <= matmult_in_a115;
    a[116] <= matmult_in_a116;
    a[117] <= matmult_in_a117;
    a[118] <= matmult_in_a118;
    a[119] <= matmult_in_a119;
    a[120] <= matmult_in_a120;
    a[121] <= matmult_in_a121;
    a[122] <= matmult_in_a122;
    a[123] <= matmult_in_a123;
    a[124] <= matmult_in_a124;
    a[125] <= matmult_in_a125;
    a[126] <= matmult_in_a126;
    a[127] <= matmult_in_a127;
    a[128] <= matmult_in_a128;
    a[129] <= matmult_in_a129;
    a[130] <= matmult_in_a130;
    a[131] <= matmult_in_a131;
    a[132] <= matmult_in_a132;
    a[133] <= matmult_in_a133;
    a[134] <= matmult_in_a134;
    a[135] <= matmult_in_a135;
    a[136] <= matmult_in_a136;
    a[137] <= matmult_in_a137;
    a[138] <= matmult_in_a138;
    a[139] <= matmult_in_a139;
    a[140] <= matmult_in_a140;
    a[141] <= matmult_in_a141;
    a[142] <= matmult_in_a142;
    a[143] <= matmult_in_a143;
    a[144] <= matmult_in_a144;
    a[145] <= matmult_in_a145;
    a[146] <= matmult_in_a146;
    a[147] <= matmult_in_a147;
    a[148] <= matmult_in_a148;
    a[149] <= matmult_in_a149;
    a[150] <= matmult_in_a150;
    a[151] <= matmult_in_a151;
    a[152] <= matmult_in_a152;
    a[153] <= matmult_in_a153;
    a[154] <= matmult_in_a154;
    a[155] <= matmult_in_a155;
    a[156] <= matmult_in_a156;
    a[157] <= matmult_in_a157;
    a[158] <= matmult_in_a158;
    a[159] <= matmult_in_a159;
    a[160] <= matmult_in_a160;
    a[161] <= matmult_in_a161;
    a[162] <= matmult_in_a162;
    a[163] <= matmult_in_a163;
    a[164] <= matmult_in_a164;
    a[165] <= matmult_in_a165;
    a[166] <= matmult_in_a166;
    a[167] <= matmult_in_a167;
    a[168] <= matmult_in_a168;
    a[169] <= matmult_in_a169;
    a[170] <= matmult_in_a170;
    a[171] <= matmult_in_a171;
    a[172] <= matmult_in_a172;
    a[173] <= matmult_in_a173;
    a[174] <= matmult_in_a174;
    a[175] <= matmult_in_a175;
    a[176] <= matmult_in_a176;
    a[177] <= matmult_in_a177;
    a[178] <= matmult_in_a178;
    a[179] <= matmult_in_a179;
    a[180] <= matmult_in_a180;
    a[181] <= matmult_in_a181;
    a[182] <= matmult_in_a182;
    a[183] <= matmult_in_a183;
    a[184] <= matmult_in_a184;
    a[185] <= matmult_in_a185;
    a[186] <= matmult_in_a186;
    a[187] <= matmult_in_a187;
    a[188] <= matmult_in_a188;
    a[189] <= matmult_in_a189;
    a[190] <= matmult_in_a190;
    a[191] <= matmult_in_a191;
    a[192] <= matmult_in_a192;
    a[193] <= matmult_in_a193;
    a[194] <= matmult_in_a194;
    a[195] <= matmult_in_a195;
    a[196] <= matmult_in_a196;
    a[197] <= matmult_in_a197;
    a[198] <= matmult_in_a198;
    a[199] <= matmult_in_a199;
    a[200] <= matmult_in_a200;
    a[201] <= matmult_in_a201;
    a[202] <= matmult_in_a202;
    a[203] <= matmult_in_a203;
    a[204] <= matmult_in_a204;
    a[205] <= matmult_in_a205;
    a[206] <= matmult_in_a206;
    a[207] <= matmult_in_a207;
    a[208] <= matmult_in_a208;
    a[209] <= matmult_in_a209;
    a[210] <= matmult_in_a210;
    a[211] <= matmult_in_a211;
    a[212] <= matmult_in_a212;
    a[213] <= matmult_in_a213;
    a[214] <= matmult_in_a214;
    a[215] <= matmult_in_a215;
    a[216] <= matmult_in_a216;
    a[217] <= matmult_in_a217;
    a[218] <= matmult_in_a218;
    a[219] <= matmult_in_a219;
    a[220] <= matmult_in_a220;
    a[221] <= matmult_in_a221;
    a[222] <= matmult_in_a222;
    a[223] <= matmult_in_a223;
    a[224] <= matmult_in_a224;
    a[225] <= matmult_in_a225;
    a[226] <= matmult_in_a226;
    a[227] <= matmult_in_a227;
    a[228] <= matmult_in_a228;
    a[229] <= matmult_in_a229;
    a[230] <= matmult_in_a230;
    a[231] <= matmult_in_a231;
    a[232] <= matmult_in_a232;
    a[233] <= matmult_in_a233;
    a[234] <= matmult_in_a234;
    a[235] <= matmult_in_a235;
    a[236] <= matmult_in_a236;
    a[237] <= matmult_in_a237;
    a[238] <= matmult_in_a238;
    a[239] <= matmult_in_a239;
    a[240] <= matmult_in_a240;
    a[241] <= matmult_in_a241;
    a[242] <= matmult_in_a242;
    a[243] <= matmult_in_a243;
    a[244] <= matmult_in_a244;
    a[245] <= matmult_in_a245;
    a[246] <= matmult_in_a246;
    a[247] <= matmult_in_a247;
    a[248] <= matmult_in_a248;
    a[249] <= matmult_in_a249;
    a[250] <= matmult_in_a250;
    a[251] <= matmult_in_a251;
    a[252] <= matmult_in_a252;
    a[253] <= matmult_in_a253;
    a[254] <= matmult_in_a254;
    a[255] <= matmult_in_a255;
    a[256] <= matmult_in_a256;
    a[257] <= matmult_in_a257;
    a[258] <= matmult_in_a258;
    a[259] <= matmult_in_a259;
    a[260] <= matmult_in_a260;
    a[261] <= matmult_in_a261;
    a[262] <= matmult_in_a262;
    a[263] <= matmult_in_a263;
    a[264] <= matmult_in_a264;
    a[265] <= matmult_in_a265;
    a[266] <= matmult_in_a266;
    a[267] <= matmult_in_a267;
    a[268] <= matmult_in_a268;
    a[269] <= matmult_in_a269;
    a[270] <= matmult_in_a270;
    a[271] <= matmult_in_a271;
    a[272] <= matmult_in_a272;
    a[273] <= matmult_in_a273;
    a[274] <= matmult_in_a274;
    a[275] <= matmult_in_a275;
    a[276] <= matmult_in_a276;
    a[277] <= matmult_in_a277;
    a[278] <= matmult_in_a278;
    a[279] <= matmult_in_a279;
    b[0] <= matmult_in_b0;
    b[1] <= matmult_in_b1;
    b[2] <= matmult_in_b2;
    b[3] <= matmult_in_b3;
    b[4] <= matmult_in_b4;
    b[5] <= matmult_in_b5;
    b[6] <= matmult_in_b6;
    b[7] <= matmult_in_b7;
    b[8] <= matmult_in_b8;
    b[9] <= matmult_in_b9;
    b[10] <= matmult_in_b10;
    b[11] <= matmult_in_b11;
    b[12] <= matmult_in_b12;
    b[13] <= matmult_in_b13;
    b[14] <= matmult_in_b14;
    b[15] <= matmult_in_b15;
    b[16] <= matmult_in_b16;
    b[17] <= matmult_in_b17;
    b[18] <= matmult_in_b18;
    b[19] <= matmult_in_b19;
    b[20] <= matmult_in_b20;
    b[21] <= matmult_in_b21;
    b[22] <= matmult_in_b22;
    b[23] <= matmult_in_b23;
    b[24] <= matmult_in_b24;
    b[25] <= matmult_in_b25;
    b[26] <= matmult_in_b26;
    b[27] <= matmult_in_b27;
    b[28] <= matmult_in_b28;
    b[29] <= matmult_in_b29;
    b[30] <= matmult_in_b30;
    b[31] <= matmult_in_b31;
    b[32] <= matmult_in_b32;
    b[33] <= matmult_in_b33;
    b[34] <= matmult_in_b34;
    b[35] <= matmult_in_b35;
    b[36] <= matmult_in_b36;
    b[37] <= matmult_in_b37;
    b[38] <= matmult_in_b38;
    b[39] <= matmult_in_b39;
    b[40] <= matmult_in_b40;
    b[41] <= matmult_in_b41;
    b[42] <= matmult_in_b42;
    b[43] <= matmult_in_b43;
    b[44] <= matmult_in_b44;
    b[45] <= matmult_in_b45;
    b[46] <= matmult_in_b46;
    b[47] <= matmult_in_b47;
    b[48] <= matmult_in_b48;
    b[49] <= matmult_in_b49;
    b[50] <= matmult_in_b50;
    b[51] <= matmult_in_b51;
    b[52] <= matmult_in_b52;
    b[53] <= matmult_in_b53;
    b[54] <= matmult_in_b54;
    b[55] <= matmult_in_b55;
    b[56] <= matmult_in_b56;
    b[57] <= matmult_in_b57;
    b[58] <= matmult_in_b58;
    b[59] <= matmult_in_b59;
    b[60] <= matmult_in_b60;
    b[61] <= matmult_in_b61;
    b[62] <= matmult_in_b62;
    b[63] <= matmult_in_b63;
    b[64] <= matmult_in_b64;
    b[65] <= matmult_in_b65;
    b[66] <= matmult_in_b66;
    b[67] <= matmult_in_b67;
    b[68] <= matmult_in_b68;
    b[69] <= matmult_in_b69;
    b[70] <= matmult_in_b70;
    b[71] <= matmult_in_b71;
    b[72] <= matmult_in_b72;
    b[73] <= matmult_in_b73;
    b[74] <= matmult_in_b74;
    b[75] <= matmult_in_b75;
    b[76] <= matmult_in_b76;
    b[77] <= matmult_in_b77;
    b[78] <= matmult_in_b78;
    b[79] <= matmult_in_b79;
    b[80] <= matmult_in_b80;
    b[81] <= matmult_in_b81;
    b[82] <= matmult_in_b82;
    b[83] <= matmult_in_b83;
    b[84] <= matmult_in_b84;
    b[85] <= matmult_in_b85;
    b[86] <= matmult_in_b86;
    b[87] <= matmult_in_b87;
    b[88] <= matmult_in_b88;
    b[89] <= matmult_in_b89;
    b[90] <= matmult_in_b90;
    b[91] <= matmult_in_b91;
    b[92] <= matmult_in_b92;
    b[93] <= matmult_in_b93;
    b[94] <= matmult_in_b94;
    b[95] <= matmult_in_b95;
    b[96] <= matmult_in_b96;
    b[97] <= matmult_in_b97;
    b[98] <= matmult_in_b98;
    b[99] <= matmult_in_b99;
    b[100] <= matmult_in_b100;
    b[101] <= matmult_in_b101;
    b[102] <= matmult_in_b102;
    b[103] <= matmult_in_b103;
    b[104] <= matmult_in_b104;
    b[105] <= matmult_in_b105;
    b[106] <= matmult_in_b106;
    b[107] <= matmult_in_b107;
    b[108] <= matmult_in_b108;
    b[109] <= matmult_in_b109;
    b[110] <= matmult_in_b110;
    b[111] <= matmult_in_b111;
    b[112] <= matmult_in_b112;
    b[113] <= matmult_in_b113;
    b[114] <= matmult_in_b114;
    b[115] <= matmult_in_b115;
    b[116] <= matmult_in_b116;
    b[117] <= matmult_in_b117;
    b[118] <= matmult_in_b118;
    b[119] <= matmult_in_b119;
    b[120] <= matmult_in_b120;
    b[121] <= matmult_in_b121;
    b[122] <= matmult_in_b122;
    b[123] <= matmult_in_b123;
    b[124] <= matmult_in_b124;
    b[125] <= matmult_in_b125;
    b[126] <= matmult_in_b126;
    b[127] <= matmult_in_b127;
    b[128] <= matmult_in_b128;
    b[129] <= matmult_in_b129;
    b[130] <= matmult_in_b130;
    b[131] <= matmult_in_b131;
    b[132] <= matmult_in_b132;
    b[133] <= matmult_in_b133;
    b[134] <= matmult_in_b134;
    b[135] <= matmult_in_b135;
    b[136] <= matmult_in_b136;
    b[137] <= matmult_in_b137;
    b[138] <= matmult_in_b138;
    b[139] <= matmult_in_b139;
    b[140] <= matmult_in_b140;
    b[141] <= matmult_in_b141;
    b[142] <= matmult_in_b142;
    b[143] <= matmult_in_b143;
    b[144] <= matmult_in_b144;
    b[145] <= matmult_in_b145;
    b[146] <= matmult_in_b146;
    b[147] <= matmult_in_b147;
    b[148] <= matmult_in_b148;
    b[149] <= matmult_in_b149;
    b[150] <= matmult_in_b150;
    b[151] <= matmult_in_b151;
    b[152] <= matmult_in_b152;
    b[153] <= matmult_in_b153;
    b[154] <= matmult_in_b154;
    b[155] <= matmult_in_b155;
    b[156] <= matmult_in_b156;
    b[157] <= matmult_in_b157;
    b[158] <= matmult_in_b158;
    b[159] <= matmult_in_b159;
    b[160] <= matmult_in_b160;
    b[161] <= matmult_in_b161;
    b[162] <= matmult_in_b162;
    b[163] <= matmult_in_b163;
    b[164] <= matmult_in_b164;
    b[165] <= matmult_in_b165;
    b[166] <= matmult_in_b166;
    b[167] <= matmult_in_b167;
    b[168] <= matmult_in_b168;
    b[169] <= matmult_in_b169;
    b[170] <= matmult_in_b170;
    b[171] <= matmult_in_b171;
    b[172] <= matmult_in_b172;
    b[173] <= matmult_in_b173;
    b[174] <= matmult_in_b174;
    b[175] <= matmult_in_b175;
    b[176] <= matmult_in_b176;
    b[177] <= matmult_in_b177;
    b[178] <= matmult_in_b178;
    b[179] <= matmult_in_b179;
    b[180] <= matmult_in_b180;
    b[181] <= matmult_in_b181;
    b[182] <= matmult_in_b182;
    b[183] <= matmult_in_b183;
    b[184] <= matmult_in_b184;
    b[185] <= matmult_in_b185;
    b[186] <= matmult_in_b186;
    b[187] <= matmult_in_b187;
    b[188] <= matmult_in_b188;
    b[189] <= matmult_in_b189;
    b[190] <= matmult_in_b190;
    b[191] <= matmult_in_b191;
    b[192] <= matmult_in_b192;
    b[193] <= matmult_in_b193;
    b[194] <= matmult_in_b194;
    b[195] <= matmult_in_b195;
    b[196] <= matmult_in_b196;
    b[197] <= matmult_in_b197;
    b[198] <= matmult_in_b198;
    b[199] <= matmult_in_b199;
    b[200] <= matmult_in_b200;
    b[201] <= matmult_in_b201;
    b[202] <= matmult_in_b202;
    b[203] <= matmult_in_b203;
    b[204] <= matmult_in_b204;
    b[205] <= matmult_in_b205;
    b[206] <= matmult_in_b206;
    b[207] <= matmult_in_b207;
    b[208] <= matmult_in_b208;
    b[209] <= matmult_in_b209;
    b[210] <= matmult_in_b210;
    b[211] <= matmult_in_b211;
    b[212] <= matmult_in_b212;
    b[213] <= matmult_in_b213;
    b[214] <= matmult_in_b214;
    b[215] <= matmult_in_b215;
    b[216] <= matmult_in_b216;
    b[217] <= matmult_in_b217;
    b[218] <= matmult_in_b218;
    b[219] <= matmult_in_b219;
    b[220] <= matmult_in_b220;
    b[221] <= matmult_in_b221;
    b[222] <= matmult_in_b222;
    b[223] <= matmult_in_b223;
    b[224] <= matmult_in_b224;
    b[225] <= matmult_in_b225;
    b[226] <= matmult_in_b226;
    b[227] <= matmult_in_b227;
    b[228] <= matmult_in_b228;
    b[229] <= matmult_in_b229;
    b[230] <= matmult_in_b230;
    b[231] <= matmult_in_b231;
    b[232] <= matmult_in_b232;
    b[233] <= matmult_in_b233;
    b[234] <= matmult_in_b234;
    b[235] <= matmult_in_b235;
    b[236] <= matmult_in_b236;
    b[237] <= matmult_in_b237;
    b[238] <= matmult_in_b238;
    b[239] <= matmult_in_b239;
    b[240] <= matmult_in_b240;
    b[241] <= matmult_in_b241;
    b[242] <= matmult_in_b242;
    b[243] <= matmult_in_b243;
    b[244] <= matmult_in_b244;
    b[245] <= matmult_in_b245;
    b[246] <= matmult_in_b246;
    b[247] <= matmult_in_b247;
    b[248] <= matmult_in_b248;
    b[249] <= matmult_in_b249;
    b[250] <= matmult_in_b250;
    b[251] <= matmult_in_b251;
    b[252] <= matmult_in_b252;
    b[253] <= matmult_in_b253;
    b[254] <= matmult_in_b254;
    b[255] <= matmult_in_b255;
    b[256] <= matmult_in_b256;
    b[257] <= matmult_in_b257;
    b[258] <= matmult_in_b258;
    b[259] <= matmult_in_b259;
    b[260] <= matmult_in_b260;
    b[261] <= matmult_in_b261;
    b[262] <= matmult_in_b262;
    b[263] <= matmult_in_b263;
    b[264] <= matmult_in_b264;
    b[265] <= matmult_in_b265;
    b[266] <= matmult_in_b266;
    b[267] <= matmult_in_b267;
    b[268] <= matmult_in_b268;
    b[269] <= matmult_in_b269;
    b[270] <= matmult_in_b270;
    b[271] <= matmult_in_b271;
    b[272] <= matmult_in_b272;
    b[273] <= matmult_in_b273;
    b[274] <= matmult_in_b274;
    b[275] <= matmult_in_b275;
    b[276] <= matmult_in_b276;
    b[277] <= matmult_in_b277;
    b[278] <= matmult_in_b278;
    b[279] <= matmult_in_b279;
end

                end
                fin: begin
                    matmult_valid <= 1;
                end
                calc: begin
                    c[0] <= a[0] * b[0] + a[1] * b[20] + a[2] * b[40] + a[3] * b[60] + a[4] * b[80] + a[5] * b[100] + a[6] * b[120] + a[7] * b[140] + a[8] * b[160] + a[9] * b[180] + a[10] * b[200] + a[11] * b[220] + a[12] * b[240] + a[13] * b[260] + a[14] * b[280] + a[15] * b[300] + a[16] * b[320] + a[17] * b[340] + a[18] * b[360] + a[19] * b[380];
                    c[1] <= a[0] * b[1] + a[1] * b[21] + a[2] * b[41] + a[3] * b[61] + a[4] * b[81] + a[5] * b[101] + a[6] * b[121] + a[7] * b[141] + a[8] * b[161] + a[9] * b[181] + a[10] * b[201] + a[11] * b[221] + a[12] * b[241] + a[13] * b[261] + a[14] * b[281] + a[15] * b[301] + a[16] * b[321] + a[17] * b[341] + a[18] * b[361] + a[19] * b[381];
                    c[2] <= a[0] * b[2] + a[1] * b[22] + a[2] * b[42] + a[3] * b[62] + a[4] * b[82] + a[5] * b[102] + a[6] * b[122] + a[7] * b[142] + a[8] * b[162] + a[9] * b[182] + a[10] * b[202] + a[11] * b[222] + a[12] * b[242] + a[13] * b[262] + a[14] * b[282] + a[15] * b[302] + a[16] * b[322] + a[17] * b[342] + a[18] * b[362] + a[19] * b[382];
                    c[3] <= a[0] * b[3] + a[1] * b[23] + a[2] * b[43] + a[3] * b[63] + a[4] * b[83] + a[5] * b[103] + a[6] * b[123] + a[7] * b[143] + a[8] * b[163] + a[9] * b[183] + a[10] * b[203] + a[11] * b[223] + a[12] * b[243] + a[13] * b[263] + a[14] * b[283] + a[15] * b[303] + a[16] * b[323] + a[17] * b[343] + a[18] * b[363] + a[19] * b[383];
                    c[4] <= a[0] * b[4] + a[1] * b[24] + a[2] * b[44] + a[3] * b[64] + a[4] * b[84] + a[5] * b[104] + a[6] * b[124] + a[7] * b[144] + a[8] * b[164] + a[9] * b[184] + a[10] * b[204] + a[11] * b[224] + a[12] * b[244] + a[13] * b[264] + a[14] * b[284] + a[15] * b[304] + a[16] * b[324] + a[17] * b[344] + a[18] * b[364] + a[19] * b[384];
                    c[5] <= a[0] * b[5] + a[1] * b[25] + a[2] * b[45] + a[3] * b[65] + a[4] * b[85] + a[5] * b[105] + a[6] * b[125] + a[7] * b[145] + a[8] * b[165] + a[9] * b[185] + a[10] * b[205] + a[11] * b[225] + a[12] * b[245] + a[13] * b[265] + a[14] * b[285] + a[15] * b[305] + a[16] * b[325] + a[17] * b[345] + a[18] * b[365] + a[19] * b[385];
                    c[6] <= a[0] * b[6] + a[1] * b[26] + a[2] * b[46] + a[3] * b[66] + a[4] * b[86] + a[5] * b[106] + a[6] * b[126] + a[7] * b[146] + a[8] * b[166] + a[9] * b[186] + a[10] * b[206] + a[11] * b[226] + a[12] * b[246] + a[13] * b[266] + a[14] * b[286] + a[15] * b[306] + a[16] * b[326] + a[17] * b[346] + a[18] * b[366] + a[19] * b[386];
                    c[7] <= a[0] * b[7] + a[1] * b[27] + a[2] * b[47] + a[3] * b[67] + a[4] * b[87] + a[5] * b[107] + a[6] * b[127] + a[7] * b[147] + a[8] * b[167] + a[9] * b[187] + a[10] * b[207] + a[11] * b[227] + a[12] * b[247] + a[13] * b[267] + a[14] * b[287] + a[15] * b[307] + a[16] * b[327] + a[17] * b[347] + a[18] * b[367] + a[19] * b[387];
                    c[8] <= a[0] * b[8] + a[1] * b[28] + a[2] * b[48] + a[3] * b[68] + a[4] * b[88] + a[5] * b[108] + a[6] * b[128] + a[7] * b[148] + a[8] * b[168] + a[9] * b[188] + a[10] * b[208] + a[11] * b[228] + a[12] * b[248] + a[13] * b[268] + a[14] * b[288] + a[15] * b[308] + a[16] * b[328] + a[17] * b[348] + a[18] * b[368] + a[19] * b[388];
                    c[9] <= a[0] * b[9] + a[1] * b[29] + a[2] * b[49] + a[3] * b[69] + a[4] * b[89] + a[5] * b[109] + a[6] * b[129] + a[7] * b[149] + a[8] * b[169] + a[9] * b[189] + a[10] * b[209] + a[11] * b[229] + a[12] * b[249] + a[13] * b[269] + a[14] * b[289] + a[15] * b[309] + a[16] * b[329] + a[17] * b[349] + a[18] * b[369] + a[19] * b[389];
                    c[10] <= a[0] * b[10] + a[1] * b[30] + a[2] * b[50] + a[3] * b[70] + a[4] * b[90] + a[5] * b[110] + a[6] * b[130] + a[7] * b[150] + a[8] * b[170] + a[9] * b[190] + a[10] * b[210] + a[11] * b[230] + a[12] * b[250] + a[13] * b[270] + a[14] * b[290] + a[15] * b[310] + a[16] * b[330] + a[17] * b[350] + a[18] * b[370] + a[19] * b[390];
                    c[11] <= a[0] * b[11] + a[1] * b[31] + a[2] * b[51] + a[3] * b[71] + a[4] * b[91] + a[5] * b[111] + a[6] * b[131] + a[7] * b[151] + a[8] * b[171] + a[9] * b[191] + a[10] * b[211] + a[11] * b[231] + a[12] * b[251] + a[13] * b[271] + a[14] * b[291] + a[15] * b[311] + a[16] * b[331] + a[17] * b[351] + a[18] * b[371] + a[19] * b[391];
                    c[12] <= a[0] * b[12] + a[1] * b[32] + a[2] * b[52] + a[3] * b[72] + a[4] * b[92] + a[5] * b[112] + a[6] * b[132] + a[7] * b[152] + a[8] * b[172] + a[9] * b[192] + a[10] * b[212] + a[11] * b[232] + a[12] * b[252] + a[13] * b[272] + a[14] * b[292] + a[15] * b[312] + a[16] * b[332] + a[17] * b[352] + a[18] * b[372] + a[19] * b[392];
                    c[13] <= a[0] * b[13] + a[1] * b[33] + a[2] * b[53] + a[3] * b[73] + a[4] * b[93] + a[5] * b[113] + a[6] * b[133] + a[7] * b[153] + a[8] * b[173] + a[9] * b[193] + a[10] * b[213] + a[11] * b[233] + a[12] * b[253] + a[13] * b[273] + a[14] * b[293] + a[15] * b[313] + a[16] * b[333] + a[17] * b[353] + a[18] * b[373] + a[19] * b[393];
                    c[14] <= a[0] * b[14] + a[1] * b[34] + a[2] * b[54] + a[3] * b[74] + a[4] * b[94] + a[5] * b[114] + a[6] * b[134] + a[7] * b[154] + a[8] * b[174] + a[9] * b[194] + a[10] * b[214] + a[11] * b[234] + a[12] * b[254] + a[13] * b[274] + a[14] * b[294] + a[15] * b[314] + a[16] * b[334] + a[17] * b[354] + a[18] * b[374] + a[19] * b[394];
                    c[15] <= a[0] * b[15] + a[1] * b[35] + a[2] * b[55] + a[3] * b[75] + a[4] * b[95] + a[5] * b[115] + a[6] * b[135] + a[7] * b[155] + a[8] * b[175] + a[9] * b[195] + a[10] * b[215] + a[11] * b[235] + a[12] * b[255] + a[13] * b[275] + a[14] * b[295] + a[15] * b[315] + a[16] * b[335] + a[17] * b[355] + a[18] * b[375] + a[19] * b[395];
                    c[16] <= a[0] * b[16] + a[1] * b[36] + a[2] * b[56] + a[3] * b[76] + a[4] * b[96] + a[5] * b[116] + a[6] * b[136] + a[7] * b[156] + a[8] * b[176] + a[9] * b[196] + a[10] * b[216] + a[11] * b[236] + a[12] * b[256] + a[13] * b[276] + a[14] * b[296] + a[15] * b[316] + a[16] * b[336] + a[17] * b[356] + a[18] * b[376] + a[19] * b[396];
                    c[17] <= a[0] * b[17] + a[1] * b[37] + a[2] * b[57] + a[3] * b[77] + a[4] * b[97] + a[5] * b[117] + a[6] * b[137] + a[7] * b[157] + a[8] * b[177] + a[9] * b[197] + a[10] * b[217] + a[11] * b[237] + a[12] * b[257] + a[13] * b[277] + a[14] * b[297] + a[15] * b[317] + a[16] * b[337] + a[17] * b[357] + a[18] * b[377] + a[19] * b[397];
                    c[18] <= a[0] * b[18] + a[1] * b[38] + a[2] * b[58] + a[3] * b[78] + a[4] * b[98] + a[5] * b[118] + a[6] * b[138] + a[7] * b[158] + a[8] * b[178] + a[9] * b[198] + a[10] * b[218] + a[11] * b[238] + a[12] * b[258] + a[13] * b[278] + a[14] * b[298] + a[15] * b[318] + a[16] * b[338] + a[17] * b[358] + a[18] * b[378] + a[19] * b[398];
                    c[19] <= a[0] * b[19] + a[1] * b[39] + a[2] * b[59] + a[3] * b[79] + a[4] * b[99] + a[5] * b[119] + a[6] * b[139] + a[7] * b[159] + a[8] * b[179] + a[9] * b[199] + a[10] * b[219] + a[11] * b[239] + a[12] * b[259] + a[13] * b[279] + a[14] * b[299] + a[15] * b[319] + a[16] * b[339] + a[17] * b[359] + a[18] * b[379] + a[19] * b[399];
                    c[20] <= a[20] * b[0] + a[21] * b[20] + a[22] * b[40] + a[23] * b[60] + a[24] * b[80] + a[25] * b[100] + a[26] * b[120] + a[27] * b[140] + a[28] * b[160] + a[29] * b[180] + a[30] * b[200] + a[31] * b[220] + a[32] * b[240] + a[33] * b[260] + a[34] * b[280] + a[35] * b[300] + a[36] * b[320] + a[37] * b[340] + a[38] * b[360] + a[39] * b[380];
                    c[21] <= a[20] * b[1] + a[21] * b[21] + a[22] * b[41] + a[23] * b[61] + a[24] * b[81] + a[25] * b[101] + a[26] * b[121] + a[27] * b[141] + a[28] * b[161] + a[29] * b[181] + a[30] * b[201] + a[31] * b[221] + a[32] * b[241] + a[33] * b[261] + a[34] * b[281] + a[35] * b[301] + a[36] * b[321] + a[37] * b[341] + a[38] * b[361] + a[39] * b[381];
                    c[22] <= a[20] * b[2] + a[21] * b[22] + a[22] * b[42] + a[23] * b[62] + a[24] * b[82] + a[25] * b[102] + a[26] * b[122] + a[27] * b[142] + a[28] * b[162] + a[29] * b[182] + a[30] * b[202] + a[31] * b[222] + a[32] * b[242] + a[33] * b[262] + a[34] * b[282] + a[35] * b[302] + a[36] * b[322] + a[37] * b[342] + a[38] * b[362] + a[39] * b[382];
                    c[23] <= a[20] * b[3] + a[21] * b[23] + a[22] * b[43] + a[23] * b[63] + a[24] * b[83] + a[25] * b[103] + a[26] * b[123] + a[27] * b[143] + a[28] * b[163] + a[29] * b[183] + a[30] * b[203] + a[31] * b[223] + a[32] * b[243] + a[33] * b[263] + a[34] * b[283] + a[35] * b[303] + a[36] * b[323] + a[37] * b[343] + a[38] * b[363] + a[39] * b[383];
                    c[24] <= a[20] * b[4] + a[21] * b[24] + a[22] * b[44] + a[23] * b[64] + a[24] * b[84] + a[25] * b[104] + a[26] * b[124] + a[27] * b[144] + a[28] * b[164] + a[29] * b[184] + a[30] * b[204] + a[31] * b[224] + a[32] * b[244] + a[33] * b[264] + a[34] * b[284] + a[35] * b[304] + a[36] * b[324] + a[37] * b[344] + a[38] * b[364] + a[39] * b[384];
                    c[25] <= a[20] * b[5] + a[21] * b[25] + a[22] * b[45] + a[23] * b[65] + a[24] * b[85] + a[25] * b[105] + a[26] * b[125] + a[27] * b[145] + a[28] * b[165] + a[29] * b[185] + a[30] * b[205] + a[31] * b[225] + a[32] * b[245] + a[33] * b[265] + a[34] * b[285] + a[35] * b[305] + a[36] * b[325] + a[37] * b[345] + a[38] * b[365] + a[39] * b[385];
                    c[26] <= a[20] * b[6] + a[21] * b[26] + a[22] * b[46] + a[23] * b[66] + a[24] * b[86] + a[25] * b[106] + a[26] * b[126] + a[27] * b[146] + a[28] * b[166] + a[29] * b[186] + a[30] * b[206] + a[31] * b[226] + a[32] * b[246] + a[33] * b[266] + a[34] * b[286] + a[35] * b[306] + a[36] * b[326] + a[37] * b[346] + a[38] * b[366] + a[39] * b[386];
                    c[27] <= a[20] * b[7] + a[21] * b[27] + a[22] * b[47] + a[23] * b[67] + a[24] * b[87] + a[25] * b[107] + a[26] * b[127] + a[27] * b[147] + a[28] * b[167] + a[29] * b[187] + a[30] * b[207] + a[31] * b[227] + a[32] * b[247] + a[33] * b[267] + a[34] * b[287] + a[35] * b[307] + a[36] * b[327] + a[37] * b[347] + a[38] * b[367] + a[39] * b[387];
                    c[28] <= a[20] * b[8] + a[21] * b[28] + a[22] * b[48] + a[23] * b[68] + a[24] * b[88] + a[25] * b[108] + a[26] * b[128] + a[27] * b[148] + a[28] * b[168] + a[29] * b[188] + a[30] * b[208] + a[31] * b[228] + a[32] * b[248] + a[33] * b[268] + a[34] * b[288] + a[35] * b[308] + a[36] * b[328] + a[37] * b[348] + a[38] * b[368] + a[39] * b[388];
                    c[29] <= a[20] * b[9] + a[21] * b[29] + a[22] * b[49] + a[23] * b[69] + a[24] * b[89] + a[25] * b[109] + a[26] * b[129] + a[27] * b[149] + a[28] * b[169] + a[29] * b[189] + a[30] * b[209] + a[31] * b[229] + a[32] * b[249] + a[33] * b[269] + a[34] * b[289] + a[35] * b[309] + a[36] * b[329] + a[37] * b[349] + a[38] * b[369] + a[39] * b[389];
                    c[30] <= a[20] * b[10] + a[21] * b[30] + a[22] * b[50] + a[23] * b[70] + a[24] * b[90] + a[25] * b[110] + a[26] * b[130] + a[27] * b[150] + a[28] * b[170] + a[29] * b[190] + a[30] * b[210] + a[31] * b[230] + a[32] * b[250] + a[33] * b[270] + a[34] * b[290] + a[35] * b[310] + a[36] * b[330] + a[37] * b[350] + a[38] * b[370] + a[39] * b[390];
                    c[31] <= a[20] * b[11] + a[21] * b[31] + a[22] * b[51] + a[23] * b[71] + a[24] * b[91] + a[25] * b[111] + a[26] * b[131] + a[27] * b[151] + a[28] * b[171] + a[29] * b[191] + a[30] * b[211] + a[31] * b[231] + a[32] * b[251] + a[33] * b[271] + a[34] * b[291] + a[35] * b[311] + a[36] * b[331] + a[37] * b[351] + a[38] * b[371] + a[39] * b[391];
                    c[32] <= a[20] * b[12] + a[21] * b[32] + a[22] * b[52] + a[23] * b[72] + a[24] * b[92] + a[25] * b[112] + a[26] * b[132] + a[27] * b[152] + a[28] * b[172] + a[29] * b[192] + a[30] * b[212] + a[31] * b[232] + a[32] * b[252] + a[33] * b[272] + a[34] * b[292] + a[35] * b[312] + a[36] * b[332] + a[37] * b[352] + a[38] * b[372] + a[39] * b[392];
                    c[33] <= a[20] * b[13] + a[21] * b[33] + a[22] * b[53] + a[23] * b[73] + a[24] * b[93] + a[25] * b[113] + a[26] * b[133] + a[27] * b[153] + a[28] * b[173] + a[29] * b[193] + a[30] * b[213] + a[31] * b[233] + a[32] * b[253] + a[33] * b[273] + a[34] * b[293] + a[35] * b[313] + a[36] * b[333] + a[37] * b[353] + a[38] * b[373] + a[39] * b[393];
                    c[34] <= a[20] * b[14] + a[21] * b[34] + a[22] * b[54] + a[23] * b[74] + a[24] * b[94] + a[25] * b[114] + a[26] * b[134] + a[27] * b[154] + a[28] * b[174] + a[29] * b[194] + a[30] * b[214] + a[31] * b[234] + a[32] * b[254] + a[33] * b[274] + a[34] * b[294] + a[35] * b[314] + a[36] * b[334] + a[37] * b[354] + a[38] * b[374] + a[39] * b[394];
                    c[35] <= a[20] * b[15] + a[21] * b[35] + a[22] * b[55] + a[23] * b[75] + a[24] * b[95] + a[25] * b[115] + a[26] * b[135] + a[27] * b[155] + a[28] * b[175] + a[29] * b[195] + a[30] * b[215] + a[31] * b[235] + a[32] * b[255] + a[33] * b[275] + a[34] * b[295] + a[35] * b[315] + a[36] * b[335] + a[37] * b[355] + a[38] * b[375] + a[39] * b[395];
                    c[36] <= a[20] * b[16] + a[21] * b[36] + a[22] * b[56] + a[23] * b[76] + a[24] * b[96] + a[25] * b[116] + a[26] * b[136] + a[27] * b[156] + a[28] * b[176] + a[29] * b[196] + a[30] * b[216] + a[31] * b[236] + a[32] * b[256] + a[33] * b[276] + a[34] * b[296] + a[35] * b[316] + a[36] * b[336] + a[37] * b[356] + a[38] * b[376] + a[39] * b[396];
                    c[37] <= a[20] * b[17] + a[21] * b[37] + a[22] * b[57] + a[23] * b[77] + a[24] * b[97] + a[25] * b[117] + a[26] * b[137] + a[27] * b[157] + a[28] * b[177] + a[29] * b[197] + a[30] * b[217] + a[31] * b[237] + a[32] * b[257] + a[33] * b[277] + a[34] * b[297] + a[35] * b[317] + a[36] * b[337] + a[37] * b[357] + a[38] * b[377] + a[39] * b[397];
                    c[38] <= a[20] * b[18] + a[21] * b[38] + a[22] * b[58] + a[23] * b[78] + a[24] * b[98] + a[25] * b[118] + a[26] * b[138] + a[27] * b[158] + a[28] * b[178] + a[29] * b[198] + a[30] * b[218] + a[31] * b[238] + a[32] * b[258] + a[33] * b[278] + a[34] * b[298] + a[35] * b[318] + a[36] * b[338] + a[37] * b[358] + a[38] * b[378] + a[39] * b[398];
                    c[39] <= a[20] * b[19] + a[21] * b[39] + a[22] * b[59] + a[23] * b[79] + a[24] * b[99] + a[25] * b[119] + a[26] * b[139] + a[27] * b[159] + a[28] * b[179] + a[29] * b[199] + a[30] * b[219] + a[31] * b[239] + a[32] * b[259] + a[33] * b[279] + a[34] * b[299] + a[35] * b[319] + a[36] * b[339] + a[37] * b[359] + a[38] * b[379] + a[39] * b[399];
                    c[40] <= a[40] * b[0] + a[41] * b[20] + a[42] * b[40] + a[43] * b[60] + a[44] * b[80] + a[45] * b[100] + a[46] * b[120] + a[47] * b[140] + a[48] * b[160] + a[49] * b[180] + a[50] * b[200] + a[51] * b[220] + a[52] * b[240] + a[53] * b[260] + a[54] * b[280] + a[55] * b[300] + a[56] * b[320] + a[57] * b[340] + a[58] * b[360] + a[59] * b[380];
                    c[41] <= a[40] * b[1] + a[41] * b[21] + a[42] * b[41] + a[43] * b[61] + a[44] * b[81] + a[45] * b[101] + a[46] * b[121] + a[47] * b[141] + a[48] * b[161] + a[49] * b[181] + a[50] * b[201] + a[51] * b[221] + a[52] * b[241] + a[53] * b[261] + a[54] * b[281] + a[55] * b[301] + a[56] * b[321] + a[57] * b[341] + a[58] * b[361] + a[59] * b[381];
                    c[42] <= a[40] * b[2] + a[41] * b[22] + a[42] * b[42] + a[43] * b[62] + a[44] * b[82] + a[45] * b[102] + a[46] * b[122] + a[47] * b[142] + a[48] * b[162] + a[49] * b[182] + a[50] * b[202] + a[51] * b[222] + a[52] * b[242] + a[53] * b[262] + a[54] * b[282] + a[55] * b[302] + a[56] * b[322] + a[57] * b[342] + a[58] * b[362] + a[59] * b[382];
                    c[43] <= a[40] * b[3] + a[41] * b[23] + a[42] * b[43] + a[43] * b[63] + a[44] * b[83] + a[45] * b[103] + a[46] * b[123] + a[47] * b[143] + a[48] * b[163] + a[49] * b[183] + a[50] * b[203] + a[51] * b[223] + a[52] * b[243] + a[53] * b[263] + a[54] * b[283] + a[55] * b[303] + a[56] * b[323] + a[57] * b[343] + a[58] * b[363] + a[59] * b[383];
                    c[44] <= a[40] * b[4] + a[41] * b[24] + a[42] * b[44] + a[43] * b[64] + a[44] * b[84] + a[45] * b[104] + a[46] * b[124] + a[47] * b[144] + a[48] * b[164] + a[49] * b[184] + a[50] * b[204] + a[51] * b[224] + a[52] * b[244] + a[53] * b[264] + a[54] * b[284] + a[55] * b[304] + a[56] * b[324] + a[57] * b[344] + a[58] * b[364] + a[59] * b[384];
                    c[45] <= a[40] * b[5] + a[41] * b[25] + a[42] * b[45] + a[43] * b[65] + a[44] * b[85] + a[45] * b[105] + a[46] * b[125] + a[47] * b[145] + a[48] * b[165] + a[49] * b[185] + a[50] * b[205] + a[51] * b[225] + a[52] * b[245] + a[53] * b[265] + a[54] * b[285] + a[55] * b[305] + a[56] * b[325] + a[57] * b[345] + a[58] * b[365] + a[59] * b[385];
                    c[46] <= a[40] * b[6] + a[41] * b[26] + a[42] * b[46] + a[43] * b[66] + a[44] * b[86] + a[45] * b[106] + a[46] * b[126] + a[47] * b[146] + a[48] * b[166] + a[49] * b[186] + a[50] * b[206] + a[51] * b[226] + a[52] * b[246] + a[53] * b[266] + a[54] * b[286] + a[55] * b[306] + a[56] * b[326] + a[57] * b[346] + a[58] * b[366] + a[59] * b[386];
                    c[47] <= a[40] * b[7] + a[41] * b[27] + a[42] * b[47] + a[43] * b[67] + a[44] * b[87] + a[45] * b[107] + a[46] * b[127] + a[47] * b[147] + a[48] * b[167] + a[49] * b[187] + a[50] * b[207] + a[51] * b[227] + a[52] * b[247] + a[53] * b[267] + a[54] * b[287] + a[55] * b[307] + a[56] * b[327] + a[57] * b[347] + a[58] * b[367] + a[59] * b[387];
                    c[48] <= a[40] * b[8] + a[41] * b[28] + a[42] * b[48] + a[43] * b[68] + a[44] * b[88] + a[45] * b[108] + a[46] * b[128] + a[47] * b[148] + a[48] * b[168] + a[49] * b[188] + a[50] * b[208] + a[51] * b[228] + a[52] * b[248] + a[53] * b[268] + a[54] * b[288] + a[55] * b[308] + a[56] * b[328] + a[57] * b[348] + a[58] * b[368] + a[59] * b[388];
                    c[49] <= a[40] * b[9] + a[41] * b[29] + a[42] * b[49] + a[43] * b[69] + a[44] * b[89] + a[45] * b[109] + a[46] * b[129] + a[47] * b[149] + a[48] * b[169] + a[49] * b[189] + a[50] * b[209] + a[51] * b[229] + a[52] * b[249] + a[53] * b[269] + a[54] * b[289] + a[55] * b[309] + a[56] * b[329] + a[57] * b[349] + a[58] * b[369] + a[59] * b[389];
                    c[50] <= a[40] * b[10] + a[41] * b[30] + a[42] * b[50] + a[43] * b[70] + a[44] * b[90] + a[45] * b[110] + a[46] * b[130] + a[47] * b[150] + a[48] * b[170] + a[49] * b[190] + a[50] * b[210] + a[51] * b[230] + a[52] * b[250] + a[53] * b[270] + a[54] * b[290] + a[55] * b[310] + a[56] * b[330] + a[57] * b[350] + a[58] * b[370] + a[59] * b[390];
                    c[51] <= a[40] * b[11] + a[41] * b[31] + a[42] * b[51] + a[43] * b[71] + a[44] * b[91] + a[45] * b[111] + a[46] * b[131] + a[47] * b[151] + a[48] * b[171] + a[49] * b[191] + a[50] * b[211] + a[51] * b[231] + a[52] * b[251] + a[53] * b[271] + a[54] * b[291] + a[55] * b[311] + a[56] * b[331] + a[57] * b[351] + a[58] * b[371] + a[59] * b[391];
                    c[52] <= a[40] * b[12] + a[41] * b[32] + a[42] * b[52] + a[43] * b[72] + a[44] * b[92] + a[45] * b[112] + a[46] * b[132] + a[47] * b[152] + a[48] * b[172] + a[49] * b[192] + a[50] * b[212] + a[51] * b[232] + a[52] * b[252] + a[53] * b[272] + a[54] * b[292] + a[55] * b[312] + a[56] * b[332] + a[57] * b[352] + a[58] * b[372] + a[59] * b[392];
                    c[53] <= a[40] * b[13] + a[41] * b[33] + a[42] * b[53] + a[43] * b[73] + a[44] * b[93] + a[45] * b[113] + a[46] * b[133] + a[47] * b[153] + a[48] * b[173] + a[49] * b[193] + a[50] * b[213] + a[51] * b[233] + a[52] * b[253] + a[53] * b[273] + a[54] * b[293] + a[55] * b[313] + a[56] * b[333] + a[57] * b[353] + a[58] * b[373] + a[59] * b[393];
                    c[54] <= a[40] * b[14] + a[41] * b[34] + a[42] * b[54] + a[43] * b[74] + a[44] * b[94] + a[45] * b[114] + a[46] * b[134] + a[47] * b[154] + a[48] * b[174] + a[49] * b[194] + a[50] * b[214] + a[51] * b[234] + a[52] * b[254] + a[53] * b[274] + a[54] * b[294] + a[55] * b[314] + a[56] * b[334] + a[57] * b[354] + a[58] * b[374] + a[59] * b[394];
                    c[55] <= a[40] * b[15] + a[41] * b[35] + a[42] * b[55] + a[43] * b[75] + a[44] * b[95] + a[45] * b[115] + a[46] * b[135] + a[47] * b[155] + a[48] * b[175] + a[49] * b[195] + a[50] * b[215] + a[51] * b[235] + a[52] * b[255] + a[53] * b[275] + a[54] * b[295] + a[55] * b[315] + a[56] * b[335] + a[57] * b[355] + a[58] * b[375] + a[59] * b[395];
                    c[56] <= a[40] * b[16] + a[41] * b[36] + a[42] * b[56] + a[43] * b[76] + a[44] * b[96] + a[45] * b[116] + a[46] * b[136] + a[47] * b[156] + a[48] * b[176] + a[49] * b[196] + a[50] * b[216] + a[51] * b[236] + a[52] * b[256] + a[53] * b[276] + a[54] * b[296] + a[55] * b[316] + a[56] * b[336] + a[57] * b[356] + a[58] * b[376] + a[59] * b[396];
                    c[57] <= a[40] * b[17] + a[41] * b[37] + a[42] * b[57] + a[43] * b[77] + a[44] * b[97] + a[45] * b[117] + a[46] * b[137] + a[47] * b[157] + a[48] * b[177] + a[49] * b[197] + a[50] * b[217] + a[51] * b[237] + a[52] * b[257] + a[53] * b[277] + a[54] * b[297] + a[55] * b[317] + a[56] * b[337] + a[57] * b[357] + a[58] * b[377] + a[59] * b[397];
                    c[58] <= a[40] * b[18] + a[41] * b[38] + a[42] * b[58] + a[43] * b[78] + a[44] * b[98] + a[45] * b[118] + a[46] * b[138] + a[47] * b[158] + a[48] * b[178] + a[49] * b[198] + a[50] * b[218] + a[51] * b[238] + a[52] * b[258] + a[53] * b[278] + a[54] * b[298] + a[55] * b[318] + a[56] * b[338] + a[57] * b[358] + a[58] * b[378] + a[59] * b[398];
                    c[59] <= a[40] * b[19] + a[41] * b[39] + a[42] * b[59] + a[43] * b[79] + a[44] * b[99] + a[45] * b[119] + a[46] * b[139] + a[47] * b[159] + a[48] * b[179] + a[49] * b[199] + a[50] * b[219] + a[51] * b[239] + a[52] * b[259] + a[53] * b[279] + a[54] * b[299] + a[55] * b[319] + a[56] * b[339] + a[57] * b[359] + a[58] * b[379] + a[59] * b[399];
                    c[60] <= a[60] * b[0] + a[61] * b[20] + a[62] * b[40] + a[63] * b[60] + a[64] * b[80] + a[65] * b[100] + a[66] * b[120] + a[67] * b[140] + a[68] * b[160] + a[69] * b[180] + a[70] * b[200] + a[71] * b[220] + a[72] * b[240] + a[73] * b[260] + a[74] * b[280] + a[75] * b[300] + a[76] * b[320] + a[77] * b[340] + a[78] * b[360] + a[79] * b[380];
                    c[61] <= a[60] * b[1] + a[61] * b[21] + a[62] * b[41] + a[63] * b[61] + a[64] * b[81] + a[65] * b[101] + a[66] * b[121] + a[67] * b[141] + a[68] * b[161] + a[69] * b[181] + a[70] * b[201] + a[71] * b[221] + a[72] * b[241] + a[73] * b[261] + a[74] * b[281] + a[75] * b[301] + a[76] * b[321] + a[77] * b[341] + a[78] * b[361] + a[79] * b[381];
                    c[62] <= a[60] * b[2] + a[61] * b[22] + a[62] * b[42] + a[63] * b[62] + a[64] * b[82] + a[65] * b[102] + a[66] * b[122] + a[67] * b[142] + a[68] * b[162] + a[69] * b[182] + a[70] * b[202] + a[71] * b[222] + a[72] * b[242] + a[73] * b[262] + a[74] * b[282] + a[75] * b[302] + a[76] * b[322] + a[77] * b[342] + a[78] * b[362] + a[79] * b[382];
                    c[63] <= a[60] * b[3] + a[61] * b[23] + a[62] * b[43] + a[63] * b[63] + a[64] * b[83] + a[65] * b[103] + a[66] * b[123] + a[67] * b[143] + a[68] * b[163] + a[69] * b[183] + a[70] * b[203] + a[71] * b[223] + a[72] * b[243] + a[73] * b[263] + a[74] * b[283] + a[75] * b[303] + a[76] * b[323] + a[77] * b[343] + a[78] * b[363] + a[79] * b[383];
                    c[64] <= a[60] * b[4] + a[61] * b[24] + a[62] * b[44] + a[63] * b[64] + a[64] * b[84] + a[65] * b[104] + a[66] * b[124] + a[67] * b[144] + a[68] * b[164] + a[69] * b[184] + a[70] * b[204] + a[71] * b[224] + a[72] * b[244] + a[73] * b[264] + a[74] * b[284] + a[75] * b[304] + a[76] * b[324] + a[77] * b[344] + a[78] * b[364] + a[79] * b[384];
                    c[65] <= a[60] * b[5] + a[61] * b[25] + a[62] * b[45] + a[63] * b[65] + a[64] * b[85] + a[65] * b[105] + a[66] * b[125] + a[67] * b[145] + a[68] * b[165] + a[69] * b[185] + a[70] * b[205] + a[71] * b[225] + a[72] * b[245] + a[73] * b[265] + a[74] * b[285] + a[75] * b[305] + a[76] * b[325] + a[77] * b[345] + a[78] * b[365] + a[79] * b[385];
                    c[66] <= a[60] * b[6] + a[61] * b[26] + a[62] * b[46] + a[63] * b[66] + a[64] * b[86] + a[65] * b[106] + a[66] * b[126] + a[67] * b[146] + a[68] * b[166] + a[69] * b[186] + a[70] * b[206] + a[71] * b[226] + a[72] * b[246] + a[73] * b[266] + a[74] * b[286] + a[75] * b[306] + a[76] * b[326] + a[77] * b[346] + a[78] * b[366] + a[79] * b[386];
                    c[67] <= a[60] * b[7] + a[61] * b[27] + a[62] * b[47] + a[63] * b[67] + a[64] * b[87] + a[65] * b[107] + a[66] * b[127] + a[67] * b[147] + a[68] * b[167] + a[69] * b[187] + a[70] * b[207] + a[71] * b[227] + a[72] * b[247] + a[73] * b[267] + a[74] * b[287] + a[75] * b[307] + a[76] * b[327] + a[77] * b[347] + a[78] * b[367] + a[79] * b[387];
                    c[68] <= a[60] * b[8] + a[61] * b[28] + a[62] * b[48] + a[63] * b[68] + a[64] * b[88] + a[65] * b[108] + a[66] * b[128] + a[67] * b[148] + a[68] * b[168] + a[69] * b[188] + a[70] * b[208] + a[71] * b[228] + a[72] * b[248] + a[73] * b[268] + a[74] * b[288] + a[75] * b[308] + a[76] * b[328] + a[77] * b[348] + a[78] * b[368] + a[79] * b[388];
                    c[69] <= a[60] * b[9] + a[61] * b[29] + a[62] * b[49] + a[63] * b[69] + a[64] * b[89] + a[65] * b[109] + a[66] * b[129] + a[67] * b[149] + a[68] * b[169] + a[69] * b[189] + a[70] * b[209] + a[71] * b[229] + a[72] * b[249] + a[73] * b[269] + a[74] * b[289] + a[75] * b[309] + a[76] * b[329] + a[77] * b[349] + a[78] * b[369] + a[79] * b[389];
                    c[70] <= a[60] * b[10] + a[61] * b[30] + a[62] * b[50] + a[63] * b[70] + a[64] * b[90] + a[65] * b[110] + a[66] * b[130] + a[67] * b[150] + a[68] * b[170] + a[69] * b[190] + a[70] * b[210] + a[71] * b[230] + a[72] * b[250] + a[73] * b[270] + a[74] * b[290] + a[75] * b[310] + a[76] * b[330] + a[77] * b[350] + a[78] * b[370] + a[79] * b[390];
                    c[71] <= a[60] * b[11] + a[61] * b[31] + a[62] * b[51] + a[63] * b[71] + a[64] * b[91] + a[65] * b[111] + a[66] * b[131] + a[67] * b[151] + a[68] * b[171] + a[69] * b[191] + a[70] * b[211] + a[71] * b[231] + a[72] * b[251] + a[73] * b[271] + a[74] * b[291] + a[75] * b[311] + a[76] * b[331] + a[77] * b[351] + a[78] * b[371] + a[79] * b[391];
                    c[72] <= a[60] * b[12] + a[61] * b[32] + a[62] * b[52] + a[63] * b[72] + a[64] * b[92] + a[65] * b[112] + a[66] * b[132] + a[67] * b[152] + a[68] * b[172] + a[69] * b[192] + a[70] * b[212] + a[71] * b[232] + a[72] * b[252] + a[73] * b[272] + a[74] * b[292] + a[75] * b[312] + a[76] * b[332] + a[77] * b[352] + a[78] * b[372] + a[79] * b[392];
                    c[73] <= a[60] * b[13] + a[61] * b[33] + a[62] * b[53] + a[63] * b[73] + a[64] * b[93] + a[65] * b[113] + a[66] * b[133] + a[67] * b[153] + a[68] * b[173] + a[69] * b[193] + a[70] * b[213] + a[71] * b[233] + a[72] * b[253] + a[73] * b[273] + a[74] * b[293] + a[75] * b[313] + a[76] * b[333] + a[77] * b[353] + a[78] * b[373] + a[79] * b[393];
                    c[74] <= a[60] * b[14] + a[61] * b[34] + a[62] * b[54] + a[63] * b[74] + a[64] * b[94] + a[65] * b[114] + a[66] * b[134] + a[67] * b[154] + a[68] * b[174] + a[69] * b[194] + a[70] * b[214] + a[71] * b[234] + a[72] * b[254] + a[73] * b[274] + a[74] * b[294] + a[75] * b[314] + a[76] * b[334] + a[77] * b[354] + a[78] * b[374] + a[79] * b[394];
                    c[75] <= a[60] * b[15] + a[61] * b[35] + a[62] * b[55] + a[63] * b[75] + a[64] * b[95] + a[65] * b[115] + a[66] * b[135] + a[67] * b[155] + a[68] * b[175] + a[69] * b[195] + a[70] * b[215] + a[71] * b[235] + a[72] * b[255] + a[73] * b[275] + a[74] * b[295] + a[75] * b[315] + a[76] * b[335] + a[77] * b[355] + a[78] * b[375] + a[79] * b[395];
                    c[76] <= a[60] * b[16] + a[61] * b[36] + a[62] * b[56] + a[63] * b[76] + a[64] * b[96] + a[65] * b[116] + a[66] * b[136] + a[67] * b[156] + a[68] * b[176] + a[69] * b[196] + a[70] * b[216] + a[71] * b[236] + a[72] * b[256] + a[73] * b[276] + a[74] * b[296] + a[75] * b[316] + a[76] * b[336] + a[77] * b[356] + a[78] * b[376] + a[79] * b[396];
                    c[77] <= a[60] * b[17] + a[61] * b[37] + a[62] * b[57] + a[63] * b[77] + a[64] * b[97] + a[65] * b[117] + a[66] * b[137] + a[67] * b[157] + a[68] * b[177] + a[69] * b[197] + a[70] * b[217] + a[71] * b[237] + a[72] * b[257] + a[73] * b[277] + a[74] * b[297] + a[75] * b[317] + a[76] * b[337] + a[77] * b[357] + a[78] * b[377] + a[79] * b[397];
                    c[78] <= a[60] * b[18] + a[61] * b[38] + a[62] * b[58] + a[63] * b[78] + a[64] * b[98] + a[65] * b[118] + a[66] * b[138] + a[67] * b[158] + a[68] * b[178] + a[69] * b[198] + a[70] * b[218] + a[71] * b[238] + a[72] * b[258] + a[73] * b[278] + a[74] * b[298] + a[75] * b[318] + a[76] * b[338] + a[77] * b[358] + a[78] * b[378] + a[79] * b[398];
                    c[79] <= a[60] * b[19] + a[61] * b[39] + a[62] * b[59] + a[63] * b[79] + a[64] * b[99] + a[65] * b[119] + a[66] * b[139] + a[67] * b[159] + a[68] * b[179] + a[69] * b[199] + a[70] * b[219] + a[71] * b[239] + a[72] * b[259] + a[73] * b[279] + a[74] * b[299] + a[75] * b[319] + a[76] * b[339] + a[77] * b[359] + a[78] * b[379] + a[79] * b[399];
                    c[80] <= a[80] * b[0] + a[81] * b[20] + a[82] * b[40] + a[83] * b[60] + a[84] * b[80] + a[85] * b[100] + a[86] * b[120] + a[87] * b[140] + a[88] * b[160] + a[89] * b[180] + a[90] * b[200] + a[91] * b[220] + a[92] * b[240] + a[93] * b[260] + a[94] * b[280] + a[95] * b[300] + a[96] * b[320] + a[97] * b[340] + a[98] * b[360] + a[99] * b[380];
                    c[81] <= a[80] * b[1] + a[81] * b[21] + a[82] * b[41] + a[83] * b[61] + a[84] * b[81] + a[85] * b[101] + a[86] * b[121] + a[87] * b[141] + a[88] * b[161] + a[89] * b[181] + a[90] * b[201] + a[91] * b[221] + a[92] * b[241] + a[93] * b[261] + a[94] * b[281] + a[95] * b[301] + a[96] * b[321] + a[97] * b[341] + a[98] * b[361] + a[99] * b[381];
                    c[82] <= a[80] * b[2] + a[81] * b[22] + a[82] * b[42] + a[83] * b[62] + a[84] * b[82] + a[85] * b[102] + a[86] * b[122] + a[87] * b[142] + a[88] * b[162] + a[89] * b[182] + a[90] * b[202] + a[91] * b[222] + a[92] * b[242] + a[93] * b[262] + a[94] * b[282] + a[95] * b[302] + a[96] * b[322] + a[97] * b[342] + a[98] * b[362] + a[99] * b[382];
                    c[83] <= a[80] * b[3] + a[81] * b[23] + a[82] * b[43] + a[83] * b[63] + a[84] * b[83] + a[85] * b[103] + a[86] * b[123] + a[87] * b[143] + a[88] * b[163] + a[89] * b[183] + a[90] * b[203] + a[91] * b[223] + a[92] * b[243] + a[93] * b[263] + a[94] * b[283] + a[95] * b[303] + a[96] * b[323] + a[97] * b[343] + a[98] * b[363] + a[99] * b[383];
                    c[84] <= a[80] * b[4] + a[81] * b[24] + a[82] * b[44] + a[83] * b[64] + a[84] * b[84] + a[85] * b[104] + a[86] * b[124] + a[87] * b[144] + a[88] * b[164] + a[89] * b[184] + a[90] * b[204] + a[91] * b[224] + a[92] * b[244] + a[93] * b[264] + a[94] * b[284] + a[95] * b[304] + a[96] * b[324] + a[97] * b[344] + a[98] * b[364] + a[99] * b[384];
                    c[85] <= a[80] * b[5] + a[81] * b[25] + a[82] * b[45] + a[83] * b[65] + a[84] * b[85] + a[85] * b[105] + a[86] * b[125] + a[87] * b[145] + a[88] * b[165] + a[89] * b[185] + a[90] * b[205] + a[91] * b[225] + a[92] * b[245] + a[93] * b[265] + a[94] * b[285] + a[95] * b[305] + a[96] * b[325] + a[97] * b[345] + a[98] * b[365] + a[99] * b[385];
                    c[86] <= a[80] * b[6] + a[81] * b[26] + a[82] * b[46] + a[83] * b[66] + a[84] * b[86] + a[85] * b[106] + a[86] * b[126] + a[87] * b[146] + a[88] * b[166] + a[89] * b[186] + a[90] * b[206] + a[91] * b[226] + a[92] * b[246] + a[93] * b[266] + a[94] * b[286] + a[95] * b[306] + a[96] * b[326] + a[97] * b[346] + a[98] * b[366] + a[99] * b[386];
                    c[87] <= a[80] * b[7] + a[81] * b[27] + a[82] * b[47] + a[83] * b[67] + a[84] * b[87] + a[85] * b[107] + a[86] * b[127] + a[87] * b[147] + a[88] * b[167] + a[89] * b[187] + a[90] * b[207] + a[91] * b[227] + a[92] * b[247] + a[93] * b[267] + a[94] * b[287] + a[95] * b[307] + a[96] * b[327] + a[97] * b[347] + a[98] * b[367] + a[99] * b[387];
                    c[88] <= a[80] * b[8] + a[81] * b[28] + a[82] * b[48] + a[83] * b[68] + a[84] * b[88] + a[85] * b[108] + a[86] * b[128] + a[87] * b[148] + a[88] * b[168] + a[89] * b[188] + a[90] * b[208] + a[91] * b[228] + a[92] * b[248] + a[93] * b[268] + a[94] * b[288] + a[95] * b[308] + a[96] * b[328] + a[97] * b[348] + a[98] * b[368] + a[99] * b[388];
                    c[89] <= a[80] * b[9] + a[81] * b[29] + a[82] * b[49] + a[83] * b[69] + a[84] * b[89] + a[85] * b[109] + a[86] * b[129] + a[87] * b[149] + a[88] * b[169] + a[89] * b[189] + a[90] * b[209] + a[91] * b[229] + a[92] * b[249] + a[93] * b[269] + a[94] * b[289] + a[95] * b[309] + a[96] * b[329] + a[97] * b[349] + a[98] * b[369] + a[99] * b[389];
                    c[90] <= a[80] * b[10] + a[81] * b[30] + a[82] * b[50] + a[83] * b[70] + a[84] * b[90] + a[85] * b[110] + a[86] * b[130] + a[87] * b[150] + a[88] * b[170] + a[89] * b[190] + a[90] * b[210] + a[91] * b[230] + a[92] * b[250] + a[93] * b[270] + a[94] * b[290] + a[95] * b[310] + a[96] * b[330] + a[97] * b[350] + a[98] * b[370] + a[99] * b[390];
                    c[91] <= a[80] * b[11] + a[81] * b[31] + a[82] * b[51] + a[83] * b[71] + a[84] * b[91] + a[85] * b[111] + a[86] * b[131] + a[87] * b[151] + a[88] * b[171] + a[89] * b[191] + a[90] * b[211] + a[91] * b[231] + a[92] * b[251] + a[93] * b[271] + a[94] * b[291] + a[95] * b[311] + a[96] * b[331] + a[97] * b[351] + a[98] * b[371] + a[99] * b[391];
                    c[92] <= a[80] * b[12] + a[81] * b[32] + a[82] * b[52] + a[83] * b[72] + a[84] * b[92] + a[85] * b[112] + a[86] * b[132] + a[87] * b[152] + a[88] * b[172] + a[89] * b[192] + a[90] * b[212] + a[91] * b[232] + a[92] * b[252] + a[93] * b[272] + a[94] * b[292] + a[95] * b[312] + a[96] * b[332] + a[97] * b[352] + a[98] * b[372] + a[99] * b[392];
                    c[93] <= a[80] * b[13] + a[81] * b[33] + a[82] * b[53] + a[83] * b[73] + a[84] * b[93] + a[85] * b[113] + a[86] * b[133] + a[87] * b[153] + a[88] * b[173] + a[89] * b[193] + a[90] * b[213] + a[91] * b[233] + a[92] * b[253] + a[93] * b[273] + a[94] * b[293] + a[95] * b[313] + a[96] * b[333] + a[97] * b[353] + a[98] * b[373] + a[99] * b[393];
                    c[94] <= a[80] * b[14] + a[81] * b[34] + a[82] * b[54] + a[83] * b[74] + a[84] * b[94] + a[85] * b[114] + a[86] * b[134] + a[87] * b[154] + a[88] * b[174] + a[89] * b[194] + a[90] * b[214] + a[91] * b[234] + a[92] * b[254] + a[93] * b[274] + a[94] * b[294] + a[95] * b[314] + a[96] * b[334] + a[97] * b[354] + a[98] * b[374] + a[99] * b[394];
                    c[95] <= a[80] * b[15] + a[81] * b[35] + a[82] * b[55] + a[83] * b[75] + a[84] * b[95] + a[85] * b[115] + a[86] * b[135] + a[87] * b[155] + a[88] * b[175] + a[89] * b[195] + a[90] * b[215] + a[91] * b[235] + a[92] * b[255] + a[93] * b[275] + a[94] * b[295] + a[95] * b[315] + a[96] * b[335] + a[97] * b[355] + a[98] * b[375] + a[99] * b[395];
                    c[96] <= a[80] * b[16] + a[81] * b[36] + a[82] * b[56] + a[83] * b[76] + a[84] * b[96] + a[85] * b[116] + a[86] * b[136] + a[87] * b[156] + a[88] * b[176] + a[89] * b[196] + a[90] * b[216] + a[91] * b[236] + a[92] * b[256] + a[93] * b[276] + a[94] * b[296] + a[95] * b[316] + a[96] * b[336] + a[97] * b[356] + a[98] * b[376] + a[99] * b[396];
                    c[97] <= a[80] * b[17] + a[81] * b[37] + a[82] * b[57] + a[83] * b[77] + a[84] * b[97] + a[85] * b[117] + a[86] * b[137] + a[87] * b[157] + a[88] * b[177] + a[89] * b[197] + a[90] * b[217] + a[91] * b[237] + a[92] * b[257] + a[93] * b[277] + a[94] * b[297] + a[95] * b[317] + a[96] * b[337] + a[97] * b[357] + a[98] * b[377] + a[99] * b[397];
                    c[98] <= a[80] * b[18] + a[81] * b[38] + a[82] * b[58] + a[83] * b[78] + a[84] * b[98] + a[85] * b[118] + a[86] * b[138] + a[87] * b[158] + a[88] * b[178] + a[89] * b[198] + a[90] * b[218] + a[91] * b[238] + a[92] * b[258] + a[93] * b[278] + a[94] * b[298] + a[95] * b[318] + a[96] * b[338] + a[97] * b[358] + a[98] * b[378] + a[99] * b[398];
                    c[99] <= a[80] * b[19] + a[81] * b[39] + a[82] * b[59] + a[83] * b[79] + a[84] * b[99] + a[85] * b[119] + a[86] * b[139] + a[87] * b[159] + a[88] * b[179] + a[89] * b[199] + a[90] * b[219] + a[91] * b[239] + a[92] * b[259] + a[93] * b[279] + a[94] * b[299] + a[95] * b[319] + a[96] * b[339] + a[97] * b[359] + a[98] * b[379] + a[99] * b[399];
                    c[100] <= a[100] * b[0] + a[101] * b[20] + a[102] * b[40] + a[103] * b[60] + a[104] * b[80] + a[105] * b[100] + a[106] * b[120] + a[107] * b[140] + a[108] * b[160] + a[109] * b[180] + a[110] * b[200] + a[111] * b[220] + a[112] * b[240] + a[113] * b[260] + a[114] * b[280] + a[115] * b[300] + a[116] * b[320] + a[117] * b[340] + a[118] * b[360] + a[119] * b[380];
                    c[101] <= a[100] * b[1] + a[101] * b[21] + a[102] * b[41] + a[103] * b[61] + a[104] * b[81] + a[105] * b[101] + a[106] * b[121] + a[107] * b[141] + a[108] * b[161] + a[109] * b[181] + a[110] * b[201] + a[111] * b[221] + a[112] * b[241] + a[113] * b[261] + a[114] * b[281] + a[115] * b[301] + a[116] * b[321] + a[117] * b[341] + a[118] * b[361] + a[119] * b[381];
                    c[102] <= a[100] * b[2] + a[101] * b[22] + a[102] * b[42] + a[103] * b[62] + a[104] * b[82] + a[105] * b[102] + a[106] * b[122] + a[107] * b[142] + a[108] * b[162] + a[109] * b[182] + a[110] * b[202] + a[111] * b[222] + a[112] * b[242] + a[113] * b[262] + a[114] * b[282] + a[115] * b[302] + a[116] * b[322] + a[117] * b[342] + a[118] * b[362] + a[119] * b[382];
                    c[103] <= a[100] * b[3] + a[101] * b[23] + a[102] * b[43] + a[103] * b[63] + a[104] * b[83] + a[105] * b[103] + a[106] * b[123] + a[107] * b[143] + a[108] * b[163] + a[109] * b[183] + a[110] * b[203] + a[111] * b[223] + a[112] * b[243] + a[113] * b[263] + a[114] * b[283] + a[115] * b[303] + a[116] * b[323] + a[117] * b[343] + a[118] * b[363] + a[119] * b[383];
                    c[104] <= a[100] * b[4] + a[101] * b[24] + a[102] * b[44] + a[103] * b[64] + a[104] * b[84] + a[105] * b[104] + a[106] * b[124] + a[107] * b[144] + a[108] * b[164] + a[109] * b[184] + a[110] * b[204] + a[111] * b[224] + a[112] * b[244] + a[113] * b[264] + a[114] * b[284] + a[115] * b[304] + a[116] * b[324] + a[117] * b[344] + a[118] * b[364] + a[119] * b[384];
                    c[105] <= a[100] * b[5] + a[101] * b[25] + a[102] * b[45] + a[103] * b[65] + a[104] * b[85] + a[105] * b[105] + a[106] * b[125] + a[107] * b[145] + a[108] * b[165] + a[109] * b[185] + a[110] * b[205] + a[111] * b[225] + a[112] * b[245] + a[113] * b[265] + a[114] * b[285] + a[115] * b[305] + a[116] * b[325] + a[117] * b[345] + a[118] * b[365] + a[119] * b[385];
                    c[106] <= a[100] * b[6] + a[101] * b[26] + a[102] * b[46] + a[103] * b[66] + a[104] * b[86] + a[105] * b[106] + a[106] * b[126] + a[107] * b[146] + a[108] * b[166] + a[109] * b[186] + a[110] * b[206] + a[111] * b[226] + a[112] * b[246] + a[113] * b[266] + a[114] * b[286] + a[115] * b[306] + a[116] * b[326] + a[117] * b[346] + a[118] * b[366] + a[119] * b[386];
                    c[107] <= a[100] * b[7] + a[101] * b[27] + a[102] * b[47] + a[103] * b[67] + a[104] * b[87] + a[105] * b[107] + a[106] * b[127] + a[107] * b[147] + a[108] * b[167] + a[109] * b[187] + a[110] * b[207] + a[111] * b[227] + a[112] * b[247] + a[113] * b[267] + a[114] * b[287] + a[115] * b[307] + a[116] * b[327] + a[117] * b[347] + a[118] * b[367] + a[119] * b[387];
                    c[108] <= a[100] * b[8] + a[101] * b[28] + a[102] * b[48] + a[103] * b[68] + a[104] * b[88] + a[105] * b[108] + a[106] * b[128] + a[107] * b[148] + a[108] * b[168] + a[109] * b[188] + a[110] * b[208] + a[111] * b[228] + a[112] * b[248] + a[113] * b[268] + a[114] * b[288] + a[115] * b[308] + a[116] * b[328] + a[117] * b[348] + a[118] * b[368] + a[119] * b[388];
                    c[109] <= a[100] * b[9] + a[101] * b[29] + a[102] * b[49] + a[103] * b[69] + a[104] * b[89] + a[105] * b[109] + a[106] * b[129] + a[107] * b[149] + a[108] * b[169] + a[109] * b[189] + a[110] * b[209] + a[111] * b[229] + a[112] * b[249] + a[113] * b[269] + a[114] * b[289] + a[115] * b[309] + a[116] * b[329] + a[117] * b[349] + a[118] * b[369] + a[119] * b[389];
                    c[110] <= a[100] * b[10] + a[101] * b[30] + a[102] * b[50] + a[103] * b[70] + a[104] * b[90] + a[105] * b[110] + a[106] * b[130] + a[107] * b[150] + a[108] * b[170] + a[109] * b[190] + a[110] * b[210] + a[111] * b[230] + a[112] * b[250] + a[113] * b[270] + a[114] * b[290] + a[115] * b[310] + a[116] * b[330] + a[117] * b[350] + a[118] * b[370] + a[119] * b[390];
                    c[111] <= a[100] * b[11] + a[101] * b[31] + a[102] * b[51] + a[103] * b[71] + a[104] * b[91] + a[105] * b[111] + a[106] * b[131] + a[107] * b[151] + a[108] * b[171] + a[109] * b[191] + a[110] * b[211] + a[111] * b[231] + a[112] * b[251] + a[113] * b[271] + a[114] * b[291] + a[115] * b[311] + a[116] * b[331] + a[117] * b[351] + a[118] * b[371] + a[119] * b[391];
                    c[112] <= a[100] * b[12] + a[101] * b[32] + a[102] * b[52] + a[103] * b[72] + a[104] * b[92] + a[105] * b[112] + a[106] * b[132] + a[107] * b[152] + a[108] * b[172] + a[109] * b[192] + a[110] * b[212] + a[111] * b[232] + a[112] * b[252] + a[113] * b[272] + a[114] * b[292] + a[115] * b[312] + a[116] * b[332] + a[117] * b[352] + a[118] * b[372] + a[119] * b[392];
                    c[113] <= a[100] * b[13] + a[101] * b[33] + a[102] * b[53] + a[103] * b[73] + a[104] * b[93] + a[105] * b[113] + a[106] * b[133] + a[107] * b[153] + a[108] * b[173] + a[109] * b[193] + a[110] * b[213] + a[111] * b[233] + a[112] * b[253] + a[113] * b[273] + a[114] * b[293] + a[115] * b[313] + a[116] * b[333] + a[117] * b[353] + a[118] * b[373] + a[119] * b[393];
                    c[114] <= a[100] * b[14] + a[101] * b[34] + a[102] * b[54] + a[103] * b[74] + a[104] * b[94] + a[105] * b[114] + a[106] * b[134] + a[107] * b[154] + a[108] * b[174] + a[109] * b[194] + a[110] * b[214] + a[111] * b[234] + a[112] * b[254] + a[113] * b[274] + a[114] * b[294] + a[115] * b[314] + a[116] * b[334] + a[117] * b[354] + a[118] * b[374] + a[119] * b[394];
                    c[115] <= a[100] * b[15] + a[101] * b[35] + a[102] * b[55] + a[103] * b[75] + a[104] * b[95] + a[105] * b[115] + a[106] * b[135] + a[107] * b[155] + a[108] * b[175] + a[109] * b[195] + a[110] * b[215] + a[111] * b[235] + a[112] * b[255] + a[113] * b[275] + a[114] * b[295] + a[115] * b[315] + a[116] * b[335] + a[117] * b[355] + a[118] * b[375] + a[119] * b[395];
                    c[116] <= a[100] * b[16] + a[101] * b[36] + a[102] * b[56] + a[103] * b[76] + a[104] * b[96] + a[105] * b[116] + a[106] * b[136] + a[107] * b[156] + a[108] * b[176] + a[109] * b[196] + a[110] * b[216] + a[111] * b[236] + a[112] * b[256] + a[113] * b[276] + a[114] * b[296] + a[115] * b[316] + a[116] * b[336] + a[117] * b[356] + a[118] * b[376] + a[119] * b[396];
                    c[117] <= a[100] * b[17] + a[101] * b[37] + a[102] * b[57] + a[103] * b[77] + a[104] * b[97] + a[105] * b[117] + a[106] * b[137] + a[107] * b[157] + a[108] * b[177] + a[109] * b[197] + a[110] * b[217] + a[111] * b[237] + a[112] * b[257] + a[113] * b[277] + a[114] * b[297] + a[115] * b[317] + a[116] * b[337] + a[117] * b[357] + a[118] * b[377] + a[119] * b[397];
                    c[118] <= a[100] * b[18] + a[101] * b[38] + a[102] * b[58] + a[103] * b[78] + a[104] * b[98] + a[105] * b[118] + a[106] * b[138] + a[107] * b[158] + a[108] * b[178] + a[109] * b[198] + a[110] * b[218] + a[111] * b[238] + a[112] * b[258] + a[113] * b[278] + a[114] * b[298] + a[115] * b[318] + a[116] * b[338] + a[117] * b[358] + a[118] * b[378] + a[119] * b[398];
                    c[119] <= a[100] * b[19] + a[101] * b[39] + a[102] * b[59] + a[103] * b[79] + a[104] * b[99] + a[105] * b[119] + a[106] * b[139] + a[107] * b[159] + a[108] * b[179] + a[109] * b[199] + a[110] * b[219] + a[111] * b[239] + a[112] * b[259] + a[113] * b[279] + a[114] * b[299] + a[115] * b[319] + a[116] * b[339] + a[117] * b[359] + a[118] * b[379] + a[119] * b[399];
                    c[120] <= a[120] * b[0] + a[121] * b[20] + a[122] * b[40] + a[123] * b[60] + a[124] * b[80] + a[125] * b[100] + a[126] * b[120] + a[127] * b[140] + a[128] * b[160] + a[129] * b[180] + a[130] * b[200] + a[131] * b[220] + a[132] * b[240] + a[133] * b[260] + a[134] * b[280] + a[135] * b[300] + a[136] * b[320] + a[137] * b[340] + a[138] * b[360] + a[139] * b[380];
                    c[121] <= a[120] * b[1] + a[121] * b[21] + a[122] * b[41] + a[123] * b[61] + a[124] * b[81] + a[125] * b[101] + a[126] * b[121] + a[127] * b[141] + a[128] * b[161] + a[129] * b[181] + a[130] * b[201] + a[131] * b[221] + a[132] * b[241] + a[133] * b[261] + a[134] * b[281] + a[135] * b[301] + a[136] * b[321] + a[137] * b[341] + a[138] * b[361] + a[139] * b[381];
                    c[122] <= a[120] * b[2] + a[121] * b[22] + a[122] * b[42] + a[123] * b[62] + a[124] * b[82] + a[125] * b[102] + a[126] * b[122] + a[127] * b[142] + a[128] * b[162] + a[129] * b[182] + a[130] * b[202] + a[131] * b[222] + a[132] * b[242] + a[133] * b[262] + a[134] * b[282] + a[135] * b[302] + a[136] * b[322] + a[137] * b[342] + a[138] * b[362] + a[139] * b[382];
                    c[123] <= a[120] * b[3] + a[121] * b[23] + a[122] * b[43] + a[123] * b[63] + a[124] * b[83] + a[125] * b[103] + a[126] * b[123] + a[127] * b[143] + a[128] * b[163] + a[129] * b[183] + a[130] * b[203] + a[131] * b[223] + a[132] * b[243] + a[133] * b[263] + a[134] * b[283] + a[135] * b[303] + a[136] * b[323] + a[137] * b[343] + a[138] * b[363] + a[139] * b[383];
                    c[124] <= a[120] * b[4] + a[121] * b[24] + a[122] * b[44] + a[123] * b[64] + a[124] * b[84] + a[125] * b[104] + a[126] * b[124] + a[127] * b[144] + a[128] * b[164] + a[129] * b[184] + a[130] * b[204] + a[131] * b[224] + a[132] * b[244] + a[133] * b[264] + a[134] * b[284] + a[135] * b[304] + a[136] * b[324] + a[137] * b[344] + a[138] * b[364] + a[139] * b[384];
                    c[125] <= a[120] * b[5] + a[121] * b[25] + a[122] * b[45] + a[123] * b[65] + a[124] * b[85] + a[125] * b[105] + a[126] * b[125] + a[127] * b[145] + a[128] * b[165] + a[129] * b[185] + a[130] * b[205] + a[131] * b[225] + a[132] * b[245] + a[133] * b[265] + a[134] * b[285] + a[135] * b[305] + a[136] * b[325] + a[137] * b[345] + a[138] * b[365] + a[139] * b[385];
                    c[126] <= a[120] * b[6] + a[121] * b[26] + a[122] * b[46] + a[123] * b[66] + a[124] * b[86] + a[125] * b[106] + a[126] * b[126] + a[127] * b[146] + a[128] * b[166] + a[129] * b[186] + a[130] * b[206] + a[131] * b[226] + a[132] * b[246] + a[133] * b[266] + a[134] * b[286] + a[135] * b[306] + a[136] * b[326] + a[137] * b[346] + a[138] * b[366] + a[139] * b[386];
                    c[127] <= a[120] * b[7] + a[121] * b[27] + a[122] * b[47] + a[123] * b[67] + a[124] * b[87] + a[125] * b[107] + a[126] * b[127] + a[127] * b[147] + a[128] * b[167] + a[129] * b[187] + a[130] * b[207] + a[131] * b[227] + a[132] * b[247] + a[133] * b[267] + a[134] * b[287] + a[135] * b[307] + a[136] * b[327] + a[137] * b[347] + a[138] * b[367] + a[139] * b[387];
                    c[128] <= a[120] * b[8] + a[121] * b[28] + a[122] * b[48] + a[123] * b[68] + a[124] * b[88] + a[125] * b[108] + a[126] * b[128] + a[127] * b[148] + a[128] * b[168] + a[129] * b[188] + a[130] * b[208] + a[131] * b[228] + a[132] * b[248] + a[133] * b[268] + a[134] * b[288] + a[135] * b[308] + a[136] * b[328] + a[137] * b[348] + a[138] * b[368] + a[139] * b[388];
                    c[129] <= a[120] * b[9] + a[121] * b[29] + a[122] * b[49] + a[123] * b[69] + a[124] * b[89] + a[125] * b[109] + a[126] * b[129] + a[127] * b[149] + a[128] * b[169] + a[129] * b[189] + a[130] * b[209] + a[131] * b[229] + a[132] * b[249] + a[133] * b[269] + a[134] * b[289] + a[135] * b[309] + a[136] * b[329] + a[137] * b[349] + a[138] * b[369] + a[139] * b[389];
                    c[130] <= a[120] * b[10] + a[121] * b[30] + a[122] * b[50] + a[123] * b[70] + a[124] * b[90] + a[125] * b[110] + a[126] * b[130] + a[127] * b[150] + a[128] * b[170] + a[129] * b[190] + a[130] * b[210] + a[131] * b[230] + a[132] * b[250] + a[133] * b[270] + a[134] * b[290] + a[135] * b[310] + a[136] * b[330] + a[137] * b[350] + a[138] * b[370] + a[139] * b[390];
                    c[131] <= a[120] * b[11] + a[121] * b[31] + a[122] * b[51] + a[123] * b[71] + a[124] * b[91] + a[125] * b[111] + a[126] * b[131] + a[127] * b[151] + a[128] * b[171] + a[129] * b[191] + a[130] * b[211] + a[131] * b[231] + a[132] * b[251] + a[133] * b[271] + a[134] * b[291] + a[135] * b[311] + a[136] * b[331] + a[137] * b[351] + a[138] * b[371] + a[139] * b[391];
                    c[132] <= a[120] * b[12] + a[121] * b[32] + a[122] * b[52] + a[123] * b[72] + a[124] * b[92] + a[125] * b[112] + a[126] * b[132] + a[127] * b[152] + a[128] * b[172] + a[129] * b[192] + a[130] * b[212] + a[131] * b[232] + a[132] * b[252] + a[133] * b[272] + a[134] * b[292] + a[135] * b[312] + a[136] * b[332] + a[137] * b[352] + a[138] * b[372] + a[139] * b[392];
                    c[133] <= a[120] * b[13] + a[121] * b[33] + a[122] * b[53] + a[123] * b[73] + a[124] * b[93] + a[125] * b[113] + a[126] * b[133] + a[127] * b[153] + a[128] * b[173] + a[129] * b[193] + a[130] * b[213] + a[131] * b[233] + a[132] * b[253] + a[133] * b[273] + a[134] * b[293] + a[135] * b[313] + a[136] * b[333] + a[137] * b[353] + a[138] * b[373] + a[139] * b[393];
                    c[134] <= a[120] * b[14] + a[121] * b[34] + a[122] * b[54] + a[123] * b[74] + a[124] * b[94] + a[125] * b[114] + a[126] * b[134] + a[127] * b[154] + a[128] * b[174] + a[129] * b[194] + a[130] * b[214] + a[131] * b[234] + a[132] * b[254] + a[133] * b[274] + a[134] * b[294] + a[135] * b[314] + a[136] * b[334] + a[137] * b[354] + a[138] * b[374] + a[139] * b[394];
                    c[135] <= a[120] * b[15] + a[121] * b[35] + a[122] * b[55] + a[123] * b[75] + a[124] * b[95] + a[125] * b[115] + a[126] * b[135] + a[127] * b[155] + a[128] * b[175] + a[129] * b[195] + a[130] * b[215] + a[131] * b[235] + a[132] * b[255] + a[133] * b[275] + a[134] * b[295] + a[135] * b[315] + a[136] * b[335] + a[137] * b[355] + a[138] * b[375] + a[139] * b[395];
                    c[136] <= a[120] * b[16] + a[121] * b[36] + a[122] * b[56] + a[123] * b[76] + a[124] * b[96] + a[125] * b[116] + a[126] * b[136] + a[127] * b[156] + a[128] * b[176] + a[129] * b[196] + a[130] * b[216] + a[131] * b[236] + a[132] * b[256] + a[133] * b[276] + a[134] * b[296] + a[135] * b[316] + a[136] * b[336] + a[137] * b[356] + a[138] * b[376] + a[139] * b[396];
                    c[137] <= a[120] * b[17] + a[121] * b[37] + a[122] * b[57] + a[123] * b[77] + a[124] * b[97] + a[125] * b[117] + a[126] * b[137] + a[127] * b[157] + a[128] * b[177] + a[129] * b[197] + a[130] * b[217] + a[131] * b[237] + a[132] * b[257] + a[133] * b[277] + a[134] * b[297] + a[135] * b[317] + a[136] * b[337] + a[137] * b[357] + a[138] * b[377] + a[139] * b[397];
                    c[138] <= a[120] * b[18] + a[121] * b[38] + a[122] * b[58] + a[123] * b[78] + a[124] * b[98] + a[125] * b[118] + a[126] * b[138] + a[127] * b[158] + a[128] * b[178] + a[129] * b[198] + a[130] * b[218] + a[131] * b[238] + a[132] * b[258] + a[133] * b[278] + a[134] * b[298] + a[135] * b[318] + a[136] * b[338] + a[137] * b[358] + a[138] * b[378] + a[139] * b[398];
                    c[139] <= a[120] * b[19] + a[121] * b[39] + a[122] * b[59] + a[123] * b[79] + a[124] * b[99] + a[125] * b[119] + a[126] * b[139] + a[127] * b[159] + a[128] * b[179] + a[129] * b[199] + a[130] * b[219] + a[131] * b[239] + a[132] * b[259] + a[133] * b[279] + a[134] * b[299] + a[135] * b[319] + a[136] * b[339] + a[137] * b[359] + a[138] * b[379] + a[139] * b[399];
                    c[140] <= a[140] * b[0] + a[141] * b[20] + a[142] * b[40] + a[143] * b[60] + a[144] * b[80] + a[145] * b[100] + a[146] * b[120] + a[147] * b[140] + a[148] * b[160] + a[149] * b[180] + a[150] * b[200] + a[151] * b[220] + a[152] * b[240] + a[153] * b[260] + a[154] * b[280] + a[155] * b[300] + a[156] * b[320] + a[157] * b[340] + a[158] * b[360] + a[159] * b[380];
                    c[141] <= a[140] * b[1] + a[141] * b[21] + a[142] * b[41] + a[143] * b[61] + a[144] * b[81] + a[145] * b[101] + a[146] * b[121] + a[147] * b[141] + a[148] * b[161] + a[149] * b[181] + a[150] * b[201] + a[151] * b[221] + a[152] * b[241] + a[153] * b[261] + a[154] * b[281] + a[155] * b[301] + a[156] * b[321] + a[157] * b[341] + a[158] * b[361] + a[159] * b[381];
                    c[142] <= a[140] * b[2] + a[141] * b[22] + a[142] * b[42] + a[143] * b[62] + a[144] * b[82] + a[145] * b[102] + a[146] * b[122] + a[147] * b[142] + a[148] * b[162] + a[149] * b[182] + a[150] * b[202] + a[151] * b[222] + a[152] * b[242] + a[153] * b[262] + a[154] * b[282] + a[155] * b[302] + a[156] * b[322] + a[157] * b[342] + a[158] * b[362] + a[159] * b[382];
                    c[143] <= a[140] * b[3] + a[141] * b[23] + a[142] * b[43] + a[143] * b[63] + a[144] * b[83] + a[145] * b[103] + a[146] * b[123] + a[147] * b[143] + a[148] * b[163] + a[149] * b[183] + a[150] * b[203] + a[151] * b[223] + a[152] * b[243] + a[153] * b[263] + a[154] * b[283] + a[155] * b[303] + a[156] * b[323] + a[157] * b[343] + a[158] * b[363] + a[159] * b[383];
                    c[144] <= a[140] * b[4] + a[141] * b[24] + a[142] * b[44] + a[143] * b[64] + a[144] * b[84] + a[145] * b[104] + a[146] * b[124] + a[147] * b[144] + a[148] * b[164] + a[149] * b[184] + a[150] * b[204] + a[151] * b[224] + a[152] * b[244] + a[153] * b[264] + a[154] * b[284] + a[155] * b[304] + a[156] * b[324] + a[157] * b[344] + a[158] * b[364] + a[159] * b[384];
                    c[145] <= a[140] * b[5] + a[141] * b[25] + a[142] * b[45] + a[143] * b[65] + a[144] * b[85] + a[145] * b[105] + a[146] * b[125] + a[147] * b[145] + a[148] * b[165] + a[149] * b[185] + a[150] * b[205] + a[151] * b[225] + a[152] * b[245] + a[153] * b[265] + a[154] * b[285] + a[155] * b[305] + a[156] * b[325] + a[157] * b[345] + a[158] * b[365] + a[159] * b[385];
                    c[146] <= a[140] * b[6] + a[141] * b[26] + a[142] * b[46] + a[143] * b[66] + a[144] * b[86] + a[145] * b[106] + a[146] * b[126] + a[147] * b[146] + a[148] * b[166] + a[149] * b[186] + a[150] * b[206] + a[151] * b[226] + a[152] * b[246] + a[153] * b[266] + a[154] * b[286] + a[155] * b[306] + a[156] * b[326] + a[157] * b[346] + a[158] * b[366] + a[159] * b[386];
                    c[147] <= a[140] * b[7] + a[141] * b[27] + a[142] * b[47] + a[143] * b[67] + a[144] * b[87] + a[145] * b[107] + a[146] * b[127] + a[147] * b[147] + a[148] * b[167] + a[149] * b[187] + a[150] * b[207] + a[151] * b[227] + a[152] * b[247] + a[153] * b[267] + a[154] * b[287] + a[155] * b[307] + a[156] * b[327] + a[157] * b[347] + a[158] * b[367] + a[159] * b[387];
                    c[148] <= a[140] * b[8] + a[141] * b[28] + a[142] * b[48] + a[143] * b[68] + a[144] * b[88] + a[145] * b[108] + a[146] * b[128] + a[147] * b[148] + a[148] * b[168] + a[149] * b[188] + a[150] * b[208] + a[151] * b[228] + a[152] * b[248] + a[153] * b[268] + a[154] * b[288] + a[155] * b[308] + a[156] * b[328] + a[157] * b[348] + a[158] * b[368] + a[159] * b[388];
                    c[149] <= a[140] * b[9] + a[141] * b[29] + a[142] * b[49] + a[143] * b[69] + a[144] * b[89] + a[145] * b[109] + a[146] * b[129] + a[147] * b[149] + a[148] * b[169] + a[149] * b[189] + a[150] * b[209] + a[151] * b[229] + a[152] * b[249] + a[153] * b[269] + a[154] * b[289] + a[155] * b[309] + a[156] * b[329] + a[157] * b[349] + a[158] * b[369] + a[159] * b[389];
                    c[150] <= a[140] * b[10] + a[141] * b[30] + a[142] * b[50] + a[143] * b[70] + a[144] * b[90] + a[145] * b[110] + a[146] * b[130] + a[147] * b[150] + a[148] * b[170] + a[149] * b[190] + a[150] * b[210] + a[151] * b[230] + a[152] * b[250] + a[153] * b[270] + a[154] * b[290] + a[155] * b[310] + a[156] * b[330] + a[157] * b[350] + a[158] * b[370] + a[159] * b[390];
                    c[151] <= a[140] * b[11] + a[141] * b[31] + a[142] * b[51] + a[143] * b[71] + a[144] * b[91] + a[145] * b[111] + a[146] * b[131] + a[147] * b[151] + a[148] * b[171] + a[149] * b[191] + a[150] * b[211] + a[151] * b[231] + a[152] * b[251] + a[153] * b[271] + a[154] * b[291] + a[155] * b[311] + a[156] * b[331] + a[157] * b[351] + a[158] * b[371] + a[159] * b[391];
                    c[152] <= a[140] * b[12] + a[141] * b[32] + a[142] * b[52] + a[143] * b[72] + a[144] * b[92] + a[145] * b[112] + a[146] * b[132] + a[147] * b[152] + a[148] * b[172] + a[149] * b[192] + a[150] * b[212] + a[151] * b[232] + a[152] * b[252] + a[153] * b[272] + a[154] * b[292] + a[155] * b[312] + a[156] * b[332] + a[157] * b[352] + a[158] * b[372] + a[159] * b[392];
                    c[153] <= a[140] * b[13] + a[141] * b[33] + a[142] * b[53] + a[143] * b[73] + a[144] * b[93] + a[145] * b[113] + a[146] * b[133] + a[147] * b[153] + a[148] * b[173] + a[149] * b[193] + a[150] * b[213] + a[151] * b[233] + a[152] * b[253] + a[153] * b[273] + a[154] * b[293] + a[155] * b[313] + a[156] * b[333] + a[157] * b[353] + a[158] * b[373] + a[159] * b[393];
                    c[154] <= a[140] * b[14] + a[141] * b[34] + a[142] * b[54] + a[143] * b[74] + a[144] * b[94] + a[145] * b[114] + a[146] * b[134] + a[147] * b[154] + a[148] * b[174] + a[149] * b[194] + a[150] * b[214] + a[151] * b[234] + a[152] * b[254] + a[153] * b[274] + a[154] * b[294] + a[155] * b[314] + a[156] * b[334] + a[157] * b[354] + a[158] * b[374] + a[159] * b[394];
                    c[155] <= a[140] * b[15] + a[141] * b[35] + a[142] * b[55] + a[143] * b[75] + a[144] * b[95] + a[145] * b[115] + a[146] * b[135] + a[147] * b[155] + a[148] * b[175] + a[149] * b[195] + a[150] * b[215] + a[151] * b[235] + a[152] * b[255] + a[153] * b[275] + a[154] * b[295] + a[155] * b[315] + a[156] * b[335] + a[157] * b[355] + a[158] * b[375] + a[159] * b[395];
                    c[156] <= a[140] * b[16] + a[141] * b[36] + a[142] * b[56] + a[143] * b[76] + a[144] * b[96] + a[145] * b[116] + a[146] * b[136] + a[147] * b[156] + a[148] * b[176] + a[149] * b[196] + a[150] * b[216] + a[151] * b[236] + a[152] * b[256] + a[153] * b[276] + a[154] * b[296] + a[155] * b[316] + a[156] * b[336] + a[157] * b[356] + a[158] * b[376] + a[159] * b[396];
                    c[157] <= a[140] * b[17] + a[141] * b[37] + a[142] * b[57] + a[143] * b[77] + a[144] * b[97] + a[145] * b[117] + a[146] * b[137] + a[147] * b[157] + a[148] * b[177] + a[149] * b[197] + a[150] * b[217] + a[151] * b[237] + a[152] * b[257] + a[153] * b[277] + a[154] * b[297] + a[155] * b[317] + a[156] * b[337] + a[157] * b[357] + a[158] * b[377] + a[159] * b[397];
                    c[158] <= a[140] * b[18] + a[141] * b[38] + a[142] * b[58] + a[143] * b[78] + a[144] * b[98] + a[145] * b[118] + a[146] * b[138] + a[147] * b[158] + a[148] * b[178] + a[149] * b[198] + a[150] * b[218] + a[151] * b[238] + a[152] * b[258] + a[153] * b[278] + a[154] * b[298] + a[155] * b[318] + a[156] * b[338] + a[157] * b[358] + a[158] * b[378] + a[159] * b[398];
                    c[159] <= a[140] * b[19] + a[141] * b[39] + a[142] * b[59] + a[143] * b[79] + a[144] * b[99] + a[145] * b[119] + a[146] * b[139] + a[147] * b[159] + a[148] * b[179] + a[149] * b[199] + a[150] * b[219] + a[151] * b[239] + a[152] * b[259] + a[153] * b[279] + a[154] * b[299] + a[155] * b[319] + a[156] * b[339] + a[157] * b[359] + a[158] * b[379] + a[159] * b[399];
                    c[160] <= a[160] * b[0] + a[161] * b[20] + a[162] * b[40] + a[163] * b[60] + a[164] * b[80] + a[165] * b[100] + a[166] * b[120] + a[167] * b[140] + a[168] * b[160] + a[169] * b[180] + a[170] * b[200] + a[171] * b[220] + a[172] * b[240] + a[173] * b[260] + a[174] * b[280] + a[175] * b[300] + a[176] * b[320] + a[177] * b[340] + a[178] * b[360] + a[179] * b[380];
                    c[161] <= a[160] * b[1] + a[161] * b[21] + a[162] * b[41] + a[163] * b[61] + a[164] * b[81] + a[165] * b[101] + a[166] * b[121] + a[167] * b[141] + a[168] * b[161] + a[169] * b[181] + a[170] * b[201] + a[171] * b[221] + a[172] * b[241] + a[173] * b[261] + a[174] * b[281] + a[175] * b[301] + a[176] * b[321] + a[177] * b[341] + a[178] * b[361] + a[179] * b[381];
                    c[162] <= a[160] * b[2] + a[161] * b[22] + a[162] * b[42] + a[163] * b[62] + a[164] * b[82] + a[165] * b[102] + a[166] * b[122] + a[167] * b[142] + a[168] * b[162] + a[169] * b[182] + a[170] * b[202] + a[171] * b[222] + a[172] * b[242] + a[173] * b[262] + a[174] * b[282] + a[175] * b[302] + a[176] * b[322] + a[177] * b[342] + a[178] * b[362] + a[179] * b[382];
                    c[163] <= a[160] * b[3] + a[161] * b[23] + a[162] * b[43] + a[163] * b[63] + a[164] * b[83] + a[165] * b[103] + a[166] * b[123] + a[167] * b[143] + a[168] * b[163] + a[169] * b[183] + a[170] * b[203] + a[171] * b[223] + a[172] * b[243] + a[173] * b[263] + a[174] * b[283] + a[175] * b[303] + a[176] * b[323] + a[177] * b[343] + a[178] * b[363] + a[179] * b[383];
                    c[164] <= a[160] * b[4] + a[161] * b[24] + a[162] * b[44] + a[163] * b[64] + a[164] * b[84] + a[165] * b[104] + a[166] * b[124] + a[167] * b[144] + a[168] * b[164] + a[169] * b[184] + a[170] * b[204] + a[171] * b[224] + a[172] * b[244] + a[173] * b[264] + a[174] * b[284] + a[175] * b[304] + a[176] * b[324] + a[177] * b[344] + a[178] * b[364] + a[179] * b[384];
                    c[165] <= a[160] * b[5] + a[161] * b[25] + a[162] * b[45] + a[163] * b[65] + a[164] * b[85] + a[165] * b[105] + a[166] * b[125] + a[167] * b[145] + a[168] * b[165] + a[169] * b[185] + a[170] * b[205] + a[171] * b[225] + a[172] * b[245] + a[173] * b[265] + a[174] * b[285] + a[175] * b[305] + a[176] * b[325] + a[177] * b[345] + a[178] * b[365] + a[179] * b[385];
                    c[166] <= a[160] * b[6] + a[161] * b[26] + a[162] * b[46] + a[163] * b[66] + a[164] * b[86] + a[165] * b[106] + a[166] * b[126] + a[167] * b[146] + a[168] * b[166] + a[169] * b[186] + a[170] * b[206] + a[171] * b[226] + a[172] * b[246] + a[173] * b[266] + a[174] * b[286] + a[175] * b[306] + a[176] * b[326] + a[177] * b[346] + a[178] * b[366] + a[179] * b[386];
                    c[167] <= a[160] * b[7] + a[161] * b[27] + a[162] * b[47] + a[163] * b[67] + a[164] * b[87] + a[165] * b[107] + a[166] * b[127] + a[167] * b[147] + a[168] * b[167] + a[169] * b[187] + a[170] * b[207] + a[171] * b[227] + a[172] * b[247] + a[173] * b[267] + a[174] * b[287] + a[175] * b[307] + a[176] * b[327] + a[177] * b[347] + a[178] * b[367] + a[179] * b[387];
                    c[168] <= a[160] * b[8] + a[161] * b[28] + a[162] * b[48] + a[163] * b[68] + a[164] * b[88] + a[165] * b[108] + a[166] * b[128] + a[167] * b[148] + a[168] * b[168] + a[169] * b[188] + a[170] * b[208] + a[171] * b[228] + a[172] * b[248] + a[173] * b[268] + a[174] * b[288] + a[175] * b[308] + a[176] * b[328] + a[177] * b[348] + a[178] * b[368] + a[179] * b[388];
                    c[169] <= a[160] * b[9] + a[161] * b[29] + a[162] * b[49] + a[163] * b[69] + a[164] * b[89] + a[165] * b[109] + a[166] * b[129] + a[167] * b[149] + a[168] * b[169] + a[169] * b[189] + a[170] * b[209] + a[171] * b[229] + a[172] * b[249] + a[173] * b[269] + a[174] * b[289] + a[175] * b[309] + a[176] * b[329] + a[177] * b[349] + a[178] * b[369] + a[179] * b[389];
                    c[170] <= a[160] * b[10] + a[161] * b[30] + a[162] * b[50] + a[163] * b[70] + a[164] * b[90] + a[165] * b[110] + a[166] * b[130] + a[167] * b[150] + a[168] * b[170] + a[169] * b[190] + a[170] * b[210] + a[171] * b[230] + a[172] * b[250] + a[173] * b[270] + a[174] * b[290] + a[175] * b[310] + a[176] * b[330] + a[177] * b[350] + a[178] * b[370] + a[179] * b[390];
                    c[171] <= a[160] * b[11] + a[161] * b[31] + a[162] * b[51] + a[163] * b[71] + a[164] * b[91] + a[165] * b[111] + a[166] * b[131] + a[167] * b[151] + a[168] * b[171] + a[169] * b[191] + a[170] * b[211] + a[171] * b[231] + a[172] * b[251] + a[173] * b[271] + a[174] * b[291] + a[175] * b[311] + a[176] * b[331] + a[177] * b[351] + a[178] * b[371] + a[179] * b[391];
                    c[172] <= a[160] * b[12] + a[161] * b[32] + a[162] * b[52] + a[163] * b[72] + a[164] * b[92] + a[165] * b[112] + a[166] * b[132] + a[167] * b[152] + a[168] * b[172] + a[169] * b[192] + a[170] * b[212] + a[171] * b[232] + a[172] * b[252] + a[173] * b[272] + a[174] * b[292] + a[175] * b[312] + a[176] * b[332] + a[177] * b[352] + a[178] * b[372] + a[179] * b[392];
                    c[173] <= a[160] * b[13] + a[161] * b[33] + a[162] * b[53] + a[163] * b[73] + a[164] * b[93] + a[165] * b[113] + a[166] * b[133] + a[167] * b[153] + a[168] * b[173] + a[169] * b[193] + a[170] * b[213] + a[171] * b[233] + a[172] * b[253] + a[173] * b[273] + a[174] * b[293] + a[175] * b[313] + a[176] * b[333] + a[177] * b[353] + a[178] * b[373] + a[179] * b[393];
                    c[174] <= a[160] * b[14] + a[161] * b[34] + a[162] * b[54] + a[163] * b[74] + a[164] * b[94] + a[165] * b[114] + a[166] * b[134] + a[167] * b[154] + a[168] * b[174] + a[169] * b[194] + a[170] * b[214] + a[171] * b[234] + a[172] * b[254] + a[173] * b[274] + a[174] * b[294] + a[175] * b[314] + a[176] * b[334] + a[177] * b[354] + a[178] * b[374] + a[179] * b[394];
                    c[175] <= a[160] * b[15] + a[161] * b[35] + a[162] * b[55] + a[163] * b[75] + a[164] * b[95] + a[165] * b[115] + a[166] * b[135] + a[167] * b[155] + a[168] * b[175] + a[169] * b[195] + a[170] * b[215] + a[171] * b[235] + a[172] * b[255] + a[173] * b[275] + a[174] * b[295] + a[175] * b[315] + a[176] * b[335] + a[177] * b[355] + a[178] * b[375] + a[179] * b[395];
                    c[176] <= a[160] * b[16] + a[161] * b[36] + a[162] * b[56] + a[163] * b[76] + a[164] * b[96] + a[165] * b[116] + a[166] * b[136] + a[167] * b[156] + a[168] * b[176] + a[169] * b[196] + a[170] * b[216] + a[171] * b[236] + a[172] * b[256] + a[173] * b[276] + a[174] * b[296] + a[175] * b[316] + a[176] * b[336] + a[177] * b[356] + a[178] * b[376] + a[179] * b[396];
                    c[177] <= a[160] * b[17] + a[161] * b[37] + a[162] * b[57] + a[163] * b[77] + a[164] * b[97] + a[165] * b[117] + a[166] * b[137] + a[167] * b[157] + a[168] * b[177] + a[169] * b[197] + a[170] * b[217] + a[171] * b[237] + a[172] * b[257] + a[173] * b[277] + a[174] * b[297] + a[175] * b[317] + a[176] * b[337] + a[177] * b[357] + a[178] * b[377] + a[179] * b[397];
                    c[178] <= a[160] * b[18] + a[161] * b[38] + a[162] * b[58] + a[163] * b[78] + a[164] * b[98] + a[165] * b[118] + a[166] * b[138] + a[167] * b[158] + a[168] * b[178] + a[169] * b[198] + a[170] * b[218] + a[171] * b[238] + a[172] * b[258] + a[173] * b[278] + a[174] * b[298] + a[175] * b[318] + a[176] * b[338] + a[177] * b[358] + a[178] * b[378] + a[179] * b[398];
                    c[179] <= a[160] * b[19] + a[161] * b[39] + a[162] * b[59] + a[163] * b[79] + a[164] * b[99] + a[165] * b[119] + a[166] * b[139] + a[167] * b[159] + a[168] * b[179] + a[169] * b[199] + a[170] * b[219] + a[171] * b[239] + a[172] * b[259] + a[173] * b[279] + a[174] * b[299] + a[175] * b[319] + a[176] * b[339] + a[177] * b[359] + a[178] * b[379] + a[179] * b[399];
                    c[180] <= a[180] * b[0] + a[181] * b[20] + a[182] * b[40] + a[183] * b[60] + a[184] * b[80] + a[185] * b[100] + a[186] * b[120] + a[187] * b[140] + a[188] * b[160] + a[189] * b[180] + a[190] * b[200] + a[191] * b[220] + a[192] * b[240] + a[193] * b[260] + a[194] * b[280] + a[195] * b[300] + a[196] * b[320] + a[197] * b[340] + a[198] * b[360] + a[199] * b[380];
                    c[181] <= a[180] * b[1] + a[181] * b[21] + a[182] * b[41] + a[183] * b[61] + a[184] * b[81] + a[185] * b[101] + a[186] * b[121] + a[187] * b[141] + a[188] * b[161] + a[189] * b[181] + a[190] * b[201] + a[191] * b[221] + a[192] * b[241] + a[193] * b[261] + a[194] * b[281] + a[195] * b[301] + a[196] * b[321] + a[197] * b[341] + a[198] * b[361] + a[199] * b[381];
                    c[182] <= a[180] * b[2] + a[181] * b[22] + a[182] * b[42] + a[183] * b[62] + a[184] * b[82] + a[185] * b[102] + a[186] * b[122] + a[187] * b[142] + a[188] * b[162] + a[189] * b[182] + a[190] * b[202] + a[191] * b[222] + a[192] * b[242] + a[193] * b[262] + a[194] * b[282] + a[195] * b[302] + a[196] * b[322] + a[197] * b[342] + a[198] * b[362] + a[199] * b[382];
                    c[183] <= a[180] * b[3] + a[181] * b[23] + a[182] * b[43] + a[183] * b[63] + a[184] * b[83] + a[185] * b[103] + a[186] * b[123] + a[187] * b[143] + a[188] * b[163] + a[189] * b[183] + a[190] * b[203] + a[191] * b[223] + a[192] * b[243] + a[193] * b[263] + a[194] * b[283] + a[195] * b[303] + a[196] * b[323] + a[197] * b[343] + a[198] * b[363] + a[199] * b[383];
                    c[184] <= a[180] * b[4] + a[181] * b[24] + a[182] * b[44] + a[183] * b[64] + a[184] * b[84] + a[185] * b[104] + a[186] * b[124] + a[187] * b[144] + a[188] * b[164] + a[189] * b[184] + a[190] * b[204] + a[191] * b[224] + a[192] * b[244] + a[193] * b[264] + a[194] * b[284] + a[195] * b[304] + a[196] * b[324] + a[197] * b[344] + a[198] * b[364] + a[199] * b[384];
                    c[185] <= a[180] * b[5] + a[181] * b[25] + a[182] * b[45] + a[183] * b[65] + a[184] * b[85] + a[185] * b[105] + a[186] * b[125] + a[187] * b[145] + a[188] * b[165] + a[189] * b[185] + a[190] * b[205] + a[191] * b[225] + a[192] * b[245] + a[193] * b[265] + a[194] * b[285] + a[195] * b[305] + a[196] * b[325] + a[197] * b[345] + a[198] * b[365] + a[199] * b[385];
                    c[186] <= a[180] * b[6] + a[181] * b[26] + a[182] * b[46] + a[183] * b[66] + a[184] * b[86] + a[185] * b[106] + a[186] * b[126] + a[187] * b[146] + a[188] * b[166] + a[189] * b[186] + a[190] * b[206] + a[191] * b[226] + a[192] * b[246] + a[193] * b[266] + a[194] * b[286] + a[195] * b[306] + a[196] * b[326] + a[197] * b[346] + a[198] * b[366] + a[199] * b[386];
                    c[187] <= a[180] * b[7] + a[181] * b[27] + a[182] * b[47] + a[183] * b[67] + a[184] * b[87] + a[185] * b[107] + a[186] * b[127] + a[187] * b[147] + a[188] * b[167] + a[189] * b[187] + a[190] * b[207] + a[191] * b[227] + a[192] * b[247] + a[193] * b[267] + a[194] * b[287] + a[195] * b[307] + a[196] * b[327] + a[197] * b[347] + a[198] * b[367] + a[199] * b[387];
                    c[188] <= a[180] * b[8] + a[181] * b[28] + a[182] * b[48] + a[183] * b[68] + a[184] * b[88] + a[185] * b[108] + a[186] * b[128] + a[187] * b[148] + a[188] * b[168] + a[189] * b[188] + a[190] * b[208] + a[191] * b[228] + a[192] * b[248] + a[193] * b[268] + a[194] * b[288] + a[195] * b[308] + a[196] * b[328] + a[197] * b[348] + a[198] * b[368] + a[199] * b[388];
                    c[189] <= a[180] * b[9] + a[181] * b[29] + a[182] * b[49] + a[183] * b[69] + a[184] * b[89] + a[185] * b[109] + a[186] * b[129] + a[187] * b[149] + a[188] * b[169] + a[189] * b[189] + a[190] * b[209] + a[191] * b[229] + a[192] * b[249] + a[193] * b[269] + a[194] * b[289] + a[195] * b[309] + a[196] * b[329] + a[197] * b[349] + a[198] * b[369] + a[199] * b[389];
                    c[190] <= a[180] * b[10] + a[181] * b[30] + a[182] * b[50] + a[183] * b[70] + a[184] * b[90] + a[185] * b[110] + a[186] * b[130] + a[187] * b[150] + a[188] * b[170] + a[189] * b[190] + a[190] * b[210] + a[191] * b[230] + a[192] * b[250] + a[193] * b[270] + a[194] * b[290] + a[195] * b[310] + a[196] * b[330] + a[197] * b[350] + a[198] * b[370] + a[199] * b[390];
                    c[191] <= a[180] * b[11] + a[181] * b[31] + a[182] * b[51] + a[183] * b[71] + a[184] * b[91] + a[185] * b[111] + a[186] * b[131] + a[187] * b[151] + a[188] * b[171] + a[189] * b[191] + a[190] * b[211] + a[191] * b[231] + a[192] * b[251] + a[193] * b[271] + a[194] * b[291] + a[195] * b[311] + a[196] * b[331] + a[197] * b[351] + a[198] * b[371] + a[199] * b[391];
                    c[192] <= a[180] * b[12] + a[181] * b[32] + a[182] * b[52] + a[183] * b[72] + a[184] * b[92] + a[185] * b[112] + a[186] * b[132] + a[187] * b[152] + a[188] * b[172] + a[189] * b[192] + a[190] * b[212] + a[191] * b[232] + a[192] * b[252] + a[193] * b[272] + a[194] * b[292] + a[195] * b[312] + a[196] * b[332] + a[197] * b[352] + a[198] * b[372] + a[199] * b[392];
                    c[193] <= a[180] * b[13] + a[181] * b[33] + a[182] * b[53] + a[183] * b[73] + a[184] * b[93] + a[185] * b[113] + a[186] * b[133] + a[187] * b[153] + a[188] * b[173] + a[189] * b[193] + a[190] * b[213] + a[191] * b[233] + a[192] * b[253] + a[193] * b[273] + a[194] * b[293] + a[195] * b[313] + a[196] * b[333] + a[197] * b[353] + a[198] * b[373] + a[199] * b[393];
                    c[194] <= a[180] * b[14] + a[181] * b[34] + a[182] * b[54] + a[183] * b[74] + a[184] * b[94] + a[185] * b[114] + a[186] * b[134] + a[187] * b[154] + a[188] * b[174] + a[189] * b[194] + a[190] * b[214] + a[191] * b[234] + a[192] * b[254] + a[193] * b[274] + a[194] * b[294] + a[195] * b[314] + a[196] * b[334] + a[197] * b[354] + a[198] * b[374] + a[199] * b[394];
                    c[195] <= a[180] * b[15] + a[181] * b[35] + a[182] * b[55] + a[183] * b[75] + a[184] * b[95] + a[185] * b[115] + a[186] * b[135] + a[187] * b[155] + a[188] * b[175] + a[189] * b[195] + a[190] * b[215] + a[191] * b[235] + a[192] * b[255] + a[193] * b[275] + a[194] * b[295] + a[195] * b[315] + a[196] * b[335] + a[197] * b[355] + a[198] * b[375] + a[199] * b[395];
                    c[196] <= a[180] * b[16] + a[181] * b[36] + a[182] * b[56] + a[183] * b[76] + a[184] * b[96] + a[185] * b[116] + a[186] * b[136] + a[187] * b[156] + a[188] * b[176] + a[189] * b[196] + a[190] * b[216] + a[191] * b[236] + a[192] * b[256] + a[193] * b[276] + a[194] * b[296] + a[195] * b[316] + a[196] * b[336] + a[197] * b[356] + a[198] * b[376] + a[199] * b[396];
                    c[197] <= a[180] * b[17] + a[181] * b[37] + a[182] * b[57] + a[183] * b[77] + a[184] * b[97] + a[185] * b[117] + a[186] * b[137] + a[187] * b[157] + a[188] * b[177] + a[189] * b[197] + a[190] * b[217] + a[191] * b[237] + a[192] * b[257] + a[193] * b[277] + a[194] * b[297] + a[195] * b[317] + a[196] * b[337] + a[197] * b[357] + a[198] * b[377] + a[199] * b[397];
                    c[198] <= a[180] * b[18] + a[181] * b[38] + a[182] * b[58] + a[183] * b[78] + a[184] * b[98] + a[185] * b[118] + a[186] * b[138] + a[187] * b[158] + a[188] * b[178] + a[189] * b[198] + a[190] * b[218] + a[191] * b[238] + a[192] * b[258] + a[193] * b[278] + a[194] * b[298] + a[195] * b[318] + a[196] * b[338] + a[197] * b[358] + a[198] * b[378] + a[199] * b[398];
                    c[199] <= a[180] * b[19] + a[181] * b[39] + a[182] * b[59] + a[183] * b[79] + a[184] * b[99] + a[185] * b[119] + a[186] * b[139] + a[187] * b[159] + a[188] * b[179] + a[189] * b[199] + a[190] * b[219] + a[191] * b[239] + a[192] * b[259] + a[193] * b[279] + a[194] * b[299] + a[195] * b[319] + a[196] * b[339] + a[197] * b[359] + a[198] * b[379] + a[199] * b[399];
                    c[200] <= a[200] * b[0] + a[201] * b[20] + a[202] * b[40] + a[203] * b[60] + a[204] * b[80] + a[205] * b[100] + a[206] * b[120] + a[207] * b[140] + a[208] * b[160] + a[209] * b[180] + a[210] * b[200] + a[211] * b[220] + a[212] * b[240] + a[213] * b[260] + a[214] * b[280] + a[215] * b[300] + a[216] * b[320] + a[217] * b[340] + a[218] * b[360] + a[219] * b[380];
                    c[201] <= a[200] * b[1] + a[201] * b[21] + a[202] * b[41] + a[203] * b[61] + a[204] * b[81] + a[205] * b[101] + a[206] * b[121] + a[207] * b[141] + a[208] * b[161] + a[209] * b[181] + a[210] * b[201] + a[211] * b[221] + a[212] * b[241] + a[213] * b[261] + a[214] * b[281] + a[215] * b[301] + a[216] * b[321] + a[217] * b[341] + a[218] * b[361] + a[219] * b[381];
                    c[202] <= a[200] * b[2] + a[201] * b[22] + a[202] * b[42] + a[203] * b[62] + a[204] * b[82] + a[205] * b[102] + a[206] * b[122] + a[207] * b[142] + a[208] * b[162] + a[209] * b[182] + a[210] * b[202] + a[211] * b[222] + a[212] * b[242] + a[213] * b[262] + a[214] * b[282] + a[215] * b[302] + a[216] * b[322] + a[217] * b[342] + a[218] * b[362] + a[219] * b[382];
                    c[203] <= a[200] * b[3] + a[201] * b[23] + a[202] * b[43] + a[203] * b[63] + a[204] * b[83] + a[205] * b[103] + a[206] * b[123] + a[207] * b[143] + a[208] * b[163] + a[209] * b[183] + a[210] * b[203] + a[211] * b[223] + a[212] * b[243] + a[213] * b[263] + a[214] * b[283] + a[215] * b[303] + a[216] * b[323] + a[217] * b[343] + a[218] * b[363] + a[219] * b[383];
                    c[204] <= a[200] * b[4] + a[201] * b[24] + a[202] * b[44] + a[203] * b[64] + a[204] * b[84] + a[205] * b[104] + a[206] * b[124] + a[207] * b[144] + a[208] * b[164] + a[209] * b[184] + a[210] * b[204] + a[211] * b[224] + a[212] * b[244] + a[213] * b[264] + a[214] * b[284] + a[215] * b[304] + a[216] * b[324] + a[217] * b[344] + a[218] * b[364] + a[219] * b[384];
                    c[205] <= a[200] * b[5] + a[201] * b[25] + a[202] * b[45] + a[203] * b[65] + a[204] * b[85] + a[205] * b[105] + a[206] * b[125] + a[207] * b[145] + a[208] * b[165] + a[209] * b[185] + a[210] * b[205] + a[211] * b[225] + a[212] * b[245] + a[213] * b[265] + a[214] * b[285] + a[215] * b[305] + a[216] * b[325] + a[217] * b[345] + a[218] * b[365] + a[219] * b[385];
                    c[206] <= a[200] * b[6] + a[201] * b[26] + a[202] * b[46] + a[203] * b[66] + a[204] * b[86] + a[205] * b[106] + a[206] * b[126] + a[207] * b[146] + a[208] * b[166] + a[209] * b[186] + a[210] * b[206] + a[211] * b[226] + a[212] * b[246] + a[213] * b[266] + a[214] * b[286] + a[215] * b[306] + a[216] * b[326] + a[217] * b[346] + a[218] * b[366] + a[219] * b[386];
                    c[207] <= a[200] * b[7] + a[201] * b[27] + a[202] * b[47] + a[203] * b[67] + a[204] * b[87] + a[205] * b[107] + a[206] * b[127] + a[207] * b[147] + a[208] * b[167] + a[209] * b[187] + a[210] * b[207] + a[211] * b[227] + a[212] * b[247] + a[213] * b[267] + a[214] * b[287] + a[215] * b[307] + a[216] * b[327] + a[217] * b[347] + a[218] * b[367] + a[219] * b[387];
                    c[208] <= a[200] * b[8] + a[201] * b[28] + a[202] * b[48] + a[203] * b[68] + a[204] * b[88] + a[205] * b[108] + a[206] * b[128] + a[207] * b[148] + a[208] * b[168] + a[209] * b[188] + a[210] * b[208] + a[211] * b[228] + a[212] * b[248] + a[213] * b[268] + a[214] * b[288] + a[215] * b[308] + a[216] * b[328] + a[217] * b[348] + a[218] * b[368] + a[219] * b[388];
                    c[209] <= a[200] * b[9] + a[201] * b[29] + a[202] * b[49] + a[203] * b[69] + a[204] * b[89] + a[205] * b[109] + a[206] * b[129] + a[207] * b[149] + a[208] * b[169] + a[209] * b[189] + a[210] * b[209] + a[211] * b[229] + a[212] * b[249] + a[213] * b[269] + a[214] * b[289] + a[215] * b[309] + a[216] * b[329] + a[217] * b[349] + a[218] * b[369] + a[219] * b[389];
                    c[210] <= a[200] * b[10] + a[201] * b[30] + a[202] * b[50] + a[203] * b[70] + a[204] * b[90] + a[205] * b[110] + a[206] * b[130] + a[207] * b[150] + a[208] * b[170] + a[209] * b[190] + a[210] * b[210] + a[211] * b[230] + a[212] * b[250] + a[213] * b[270] + a[214] * b[290] + a[215] * b[310] + a[216] * b[330] + a[217] * b[350] + a[218] * b[370] + a[219] * b[390];
                    c[211] <= a[200] * b[11] + a[201] * b[31] + a[202] * b[51] + a[203] * b[71] + a[204] * b[91] + a[205] * b[111] + a[206] * b[131] + a[207] * b[151] + a[208] * b[171] + a[209] * b[191] + a[210] * b[211] + a[211] * b[231] + a[212] * b[251] + a[213] * b[271] + a[214] * b[291] + a[215] * b[311] + a[216] * b[331] + a[217] * b[351] + a[218] * b[371] + a[219] * b[391];
                    c[212] <= a[200] * b[12] + a[201] * b[32] + a[202] * b[52] + a[203] * b[72] + a[204] * b[92] + a[205] * b[112] + a[206] * b[132] + a[207] * b[152] + a[208] * b[172] + a[209] * b[192] + a[210] * b[212] + a[211] * b[232] + a[212] * b[252] + a[213] * b[272] + a[214] * b[292] + a[215] * b[312] + a[216] * b[332] + a[217] * b[352] + a[218] * b[372] + a[219] * b[392];
                    c[213] <= a[200] * b[13] + a[201] * b[33] + a[202] * b[53] + a[203] * b[73] + a[204] * b[93] + a[205] * b[113] + a[206] * b[133] + a[207] * b[153] + a[208] * b[173] + a[209] * b[193] + a[210] * b[213] + a[211] * b[233] + a[212] * b[253] + a[213] * b[273] + a[214] * b[293] + a[215] * b[313] + a[216] * b[333] + a[217] * b[353] + a[218] * b[373] + a[219] * b[393];
                    c[214] <= a[200] * b[14] + a[201] * b[34] + a[202] * b[54] + a[203] * b[74] + a[204] * b[94] + a[205] * b[114] + a[206] * b[134] + a[207] * b[154] + a[208] * b[174] + a[209] * b[194] + a[210] * b[214] + a[211] * b[234] + a[212] * b[254] + a[213] * b[274] + a[214] * b[294] + a[215] * b[314] + a[216] * b[334] + a[217] * b[354] + a[218] * b[374] + a[219] * b[394];
                    c[215] <= a[200] * b[15] + a[201] * b[35] + a[202] * b[55] + a[203] * b[75] + a[204] * b[95] + a[205] * b[115] + a[206] * b[135] + a[207] * b[155] + a[208] * b[175] + a[209] * b[195] + a[210] * b[215] + a[211] * b[235] + a[212] * b[255] + a[213] * b[275] + a[214] * b[295] + a[215] * b[315] + a[216] * b[335] + a[217] * b[355] + a[218] * b[375] + a[219] * b[395];
                    c[216] <= a[200] * b[16] + a[201] * b[36] + a[202] * b[56] + a[203] * b[76] + a[204] * b[96] + a[205] * b[116] + a[206] * b[136] + a[207] * b[156] + a[208] * b[176] + a[209] * b[196] + a[210] * b[216] + a[211] * b[236] + a[212] * b[256] + a[213] * b[276] + a[214] * b[296] + a[215] * b[316] + a[216] * b[336] + a[217] * b[356] + a[218] * b[376] + a[219] * b[396];
                    c[217] <= a[200] * b[17] + a[201] * b[37] + a[202] * b[57] + a[203] * b[77] + a[204] * b[97] + a[205] * b[117] + a[206] * b[137] + a[207] * b[157] + a[208] * b[177] + a[209] * b[197] + a[210] * b[217] + a[211] * b[237] + a[212] * b[257] + a[213] * b[277] + a[214] * b[297] + a[215] * b[317] + a[216] * b[337] + a[217] * b[357] + a[218] * b[377] + a[219] * b[397];
                    c[218] <= a[200] * b[18] + a[201] * b[38] + a[202] * b[58] + a[203] * b[78] + a[204] * b[98] + a[205] * b[118] + a[206] * b[138] + a[207] * b[158] + a[208] * b[178] + a[209] * b[198] + a[210] * b[218] + a[211] * b[238] + a[212] * b[258] + a[213] * b[278] + a[214] * b[298] + a[215] * b[318] + a[216] * b[338] + a[217] * b[358] + a[218] * b[378] + a[219] * b[398];
                    c[219] <= a[200] * b[19] + a[201] * b[39] + a[202] * b[59] + a[203] * b[79] + a[204] * b[99] + a[205] * b[119] + a[206] * b[139] + a[207] * b[159] + a[208] * b[179] + a[209] * b[199] + a[210] * b[219] + a[211] * b[239] + a[212] * b[259] + a[213] * b[279] + a[214] * b[299] + a[215] * b[319] + a[216] * b[339] + a[217] * b[359] + a[218] * b[379] + a[219] * b[399];
                    c[220] <= a[220] * b[0] + a[221] * b[20] + a[222] * b[40] + a[223] * b[60] + a[224] * b[80] + a[225] * b[100] + a[226] * b[120] + a[227] * b[140] + a[228] * b[160] + a[229] * b[180] + a[230] * b[200] + a[231] * b[220] + a[232] * b[240] + a[233] * b[260] + a[234] * b[280] + a[235] * b[300] + a[236] * b[320] + a[237] * b[340] + a[238] * b[360] + a[239] * b[380];
                    c[221] <= a[220] * b[1] + a[221] * b[21] + a[222] * b[41] + a[223] * b[61] + a[224] * b[81] + a[225] * b[101] + a[226] * b[121] + a[227] * b[141] + a[228] * b[161] + a[229] * b[181] + a[230] * b[201] + a[231] * b[221] + a[232] * b[241] + a[233] * b[261] + a[234] * b[281] + a[235] * b[301] + a[236] * b[321] + a[237] * b[341] + a[238] * b[361] + a[239] * b[381];
                    c[222] <= a[220] * b[2] + a[221] * b[22] + a[222] * b[42] + a[223] * b[62] + a[224] * b[82] + a[225] * b[102] + a[226] * b[122] + a[227] * b[142] + a[228] * b[162] + a[229] * b[182] + a[230] * b[202] + a[231] * b[222] + a[232] * b[242] + a[233] * b[262] + a[234] * b[282] + a[235] * b[302] + a[236] * b[322] + a[237] * b[342] + a[238] * b[362] + a[239] * b[382];
                    c[223] <= a[220] * b[3] + a[221] * b[23] + a[222] * b[43] + a[223] * b[63] + a[224] * b[83] + a[225] * b[103] + a[226] * b[123] + a[227] * b[143] + a[228] * b[163] + a[229] * b[183] + a[230] * b[203] + a[231] * b[223] + a[232] * b[243] + a[233] * b[263] + a[234] * b[283] + a[235] * b[303] + a[236] * b[323] + a[237] * b[343] + a[238] * b[363] + a[239] * b[383];
                    c[224] <= a[220] * b[4] + a[221] * b[24] + a[222] * b[44] + a[223] * b[64] + a[224] * b[84] + a[225] * b[104] + a[226] * b[124] + a[227] * b[144] + a[228] * b[164] + a[229] * b[184] + a[230] * b[204] + a[231] * b[224] + a[232] * b[244] + a[233] * b[264] + a[234] * b[284] + a[235] * b[304] + a[236] * b[324] + a[237] * b[344] + a[238] * b[364] + a[239] * b[384];
                    c[225] <= a[220] * b[5] + a[221] * b[25] + a[222] * b[45] + a[223] * b[65] + a[224] * b[85] + a[225] * b[105] + a[226] * b[125] + a[227] * b[145] + a[228] * b[165] + a[229] * b[185] + a[230] * b[205] + a[231] * b[225] + a[232] * b[245] + a[233] * b[265] + a[234] * b[285] + a[235] * b[305] + a[236] * b[325] + a[237] * b[345] + a[238] * b[365] + a[239] * b[385];
                    c[226] <= a[220] * b[6] + a[221] * b[26] + a[222] * b[46] + a[223] * b[66] + a[224] * b[86] + a[225] * b[106] + a[226] * b[126] + a[227] * b[146] + a[228] * b[166] + a[229] * b[186] + a[230] * b[206] + a[231] * b[226] + a[232] * b[246] + a[233] * b[266] + a[234] * b[286] + a[235] * b[306] + a[236] * b[326] + a[237] * b[346] + a[238] * b[366] + a[239] * b[386];
                    c[227] <= a[220] * b[7] + a[221] * b[27] + a[222] * b[47] + a[223] * b[67] + a[224] * b[87] + a[225] * b[107] + a[226] * b[127] + a[227] * b[147] + a[228] * b[167] + a[229] * b[187] + a[230] * b[207] + a[231] * b[227] + a[232] * b[247] + a[233] * b[267] + a[234] * b[287] + a[235] * b[307] + a[236] * b[327] + a[237] * b[347] + a[238] * b[367] + a[239] * b[387];
                    c[228] <= a[220] * b[8] + a[221] * b[28] + a[222] * b[48] + a[223] * b[68] + a[224] * b[88] + a[225] * b[108] + a[226] * b[128] + a[227] * b[148] + a[228] * b[168] + a[229] * b[188] + a[230] * b[208] + a[231] * b[228] + a[232] * b[248] + a[233] * b[268] + a[234] * b[288] + a[235] * b[308] + a[236] * b[328] + a[237] * b[348] + a[238] * b[368] + a[239] * b[388];
                    c[229] <= a[220] * b[9] + a[221] * b[29] + a[222] * b[49] + a[223] * b[69] + a[224] * b[89] + a[225] * b[109] + a[226] * b[129] + a[227] * b[149] + a[228] * b[169] + a[229] * b[189] + a[230] * b[209] + a[231] * b[229] + a[232] * b[249] + a[233] * b[269] + a[234] * b[289] + a[235] * b[309] + a[236] * b[329] + a[237] * b[349] + a[238] * b[369] + a[239] * b[389];
                    c[230] <= a[220] * b[10] + a[221] * b[30] + a[222] * b[50] + a[223] * b[70] + a[224] * b[90] + a[225] * b[110] + a[226] * b[130] + a[227] * b[150] + a[228] * b[170] + a[229] * b[190] + a[230] * b[210] + a[231] * b[230] + a[232] * b[250] + a[233] * b[270] + a[234] * b[290] + a[235] * b[310] + a[236] * b[330] + a[237] * b[350] + a[238] * b[370] + a[239] * b[390];
                    c[231] <= a[220] * b[11] + a[221] * b[31] + a[222] * b[51] + a[223] * b[71] + a[224] * b[91] + a[225] * b[111] + a[226] * b[131] + a[227] * b[151] + a[228] * b[171] + a[229] * b[191] + a[230] * b[211] + a[231] * b[231] + a[232] * b[251] + a[233] * b[271] + a[234] * b[291] + a[235] * b[311] + a[236] * b[331] + a[237] * b[351] + a[238] * b[371] + a[239] * b[391];
                    c[232] <= a[220] * b[12] + a[221] * b[32] + a[222] * b[52] + a[223] * b[72] + a[224] * b[92] + a[225] * b[112] + a[226] * b[132] + a[227] * b[152] + a[228] * b[172] + a[229] * b[192] + a[230] * b[212] + a[231] * b[232] + a[232] * b[252] + a[233] * b[272] + a[234] * b[292] + a[235] * b[312] + a[236] * b[332] + a[237] * b[352] + a[238] * b[372] + a[239] * b[392];
                    c[233] <= a[220] * b[13] + a[221] * b[33] + a[222] * b[53] + a[223] * b[73] + a[224] * b[93] + a[225] * b[113] + a[226] * b[133] + a[227] * b[153] + a[228] * b[173] + a[229] * b[193] + a[230] * b[213] + a[231] * b[233] + a[232] * b[253] + a[233] * b[273] + a[234] * b[293] + a[235] * b[313] + a[236] * b[333] + a[237] * b[353] + a[238] * b[373] + a[239] * b[393];
                    c[234] <= a[220] * b[14] + a[221] * b[34] + a[222] * b[54] + a[223] * b[74] + a[224] * b[94] + a[225] * b[114] + a[226] * b[134] + a[227] * b[154] + a[228] * b[174] + a[229] * b[194] + a[230] * b[214] + a[231] * b[234] + a[232] * b[254] + a[233] * b[274] + a[234] * b[294] + a[235] * b[314] + a[236] * b[334] + a[237] * b[354] + a[238] * b[374] + a[239] * b[394];
                    c[235] <= a[220] * b[15] + a[221] * b[35] + a[222] * b[55] + a[223] * b[75] + a[224] * b[95] + a[225] * b[115] + a[226] * b[135] + a[227] * b[155] + a[228] * b[175] + a[229] * b[195] + a[230] * b[215] + a[231] * b[235] + a[232] * b[255] + a[233] * b[275] + a[234] * b[295] + a[235] * b[315] + a[236] * b[335] + a[237] * b[355] + a[238] * b[375] + a[239] * b[395];
                    c[236] <= a[220] * b[16] + a[221] * b[36] + a[222] * b[56] + a[223] * b[76] + a[224] * b[96] + a[225] * b[116] + a[226] * b[136] + a[227] * b[156] + a[228] * b[176] + a[229] * b[196] + a[230] * b[216] + a[231] * b[236] + a[232] * b[256] + a[233] * b[276] + a[234] * b[296] + a[235] * b[316] + a[236] * b[336] + a[237] * b[356] + a[238] * b[376] + a[239] * b[396];
                    c[237] <= a[220] * b[17] + a[221] * b[37] + a[222] * b[57] + a[223] * b[77] + a[224] * b[97] + a[225] * b[117] + a[226] * b[137] + a[227] * b[157] + a[228] * b[177] + a[229] * b[197] + a[230] * b[217] + a[231] * b[237] + a[232] * b[257] + a[233] * b[277] + a[234] * b[297] + a[235] * b[317] + a[236] * b[337] + a[237] * b[357] + a[238] * b[377] + a[239] * b[397];
                    c[238] <= a[220] * b[18] + a[221] * b[38] + a[222] * b[58] + a[223] * b[78] + a[224] * b[98] + a[225] * b[118] + a[226] * b[138] + a[227] * b[158] + a[228] * b[178] + a[229] * b[198] + a[230] * b[218] + a[231] * b[238] + a[232] * b[258] + a[233] * b[278] + a[234] * b[298] + a[235] * b[318] + a[236] * b[338] + a[237] * b[358] + a[238] * b[378] + a[239] * b[398];
                    c[239] <= a[220] * b[19] + a[221] * b[39] + a[222] * b[59] + a[223] * b[79] + a[224] * b[99] + a[225] * b[119] + a[226] * b[139] + a[227] * b[159] + a[228] * b[179] + a[229] * b[199] + a[230] * b[219] + a[231] * b[239] + a[232] * b[259] + a[233] * b[279] + a[234] * b[299] + a[235] * b[319] + a[236] * b[339] + a[237] * b[359] + a[238] * b[379] + a[239] * b[399];
                    c[240] <= a[240] * b[0] + a[241] * b[20] + a[242] * b[40] + a[243] * b[60] + a[244] * b[80] + a[245] * b[100] + a[246] * b[120] + a[247] * b[140] + a[248] * b[160] + a[249] * b[180] + a[250] * b[200] + a[251] * b[220] + a[252] * b[240] + a[253] * b[260] + a[254] * b[280] + a[255] * b[300] + a[256] * b[320] + a[257] * b[340] + a[258] * b[360] + a[259] * b[380];
                    c[241] <= a[240] * b[1] + a[241] * b[21] + a[242] * b[41] + a[243] * b[61] + a[244] * b[81] + a[245] * b[101] + a[246] * b[121] + a[247] * b[141] + a[248] * b[161] + a[249] * b[181] + a[250] * b[201] + a[251] * b[221] + a[252] * b[241] + a[253] * b[261] + a[254] * b[281] + a[255] * b[301] + a[256] * b[321] + a[257] * b[341] + a[258] * b[361] + a[259] * b[381];
                    c[242] <= a[240] * b[2] + a[241] * b[22] + a[242] * b[42] + a[243] * b[62] + a[244] * b[82] + a[245] * b[102] + a[246] * b[122] + a[247] * b[142] + a[248] * b[162] + a[249] * b[182] + a[250] * b[202] + a[251] * b[222] + a[252] * b[242] + a[253] * b[262] + a[254] * b[282] + a[255] * b[302] + a[256] * b[322] + a[257] * b[342] + a[258] * b[362] + a[259] * b[382];
                    c[243] <= a[240] * b[3] + a[241] * b[23] + a[242] * b[43] + a[243] * b[63] + a[244] * b[83] + a[245] * b[103] + a[246] * b[123] + a[247] * b[143] + a[248] * b[163] + a[249] * b[183] + a[250] * b[203] + a[251] * b[223] + a[252] * b[243] + a[253] * b[263] + a[254] * b[283] + a[255] * b[303] + a[256] * b[323] + a[257] * b[343] + a[258] * b[363] + a[259] * b[383];
                    c[244] <= a[240] * b[4] + a[241] * b[24] + a[242] * b[44] + a[243] * b[64] + a[244] * b[84] + a[245] * b[104] + a[246] * b[124] + a[247] * b[144] + a[248] * b[164] + a[249] * b[184] + a[250] * b[204] + a[251] * b[224] + a[252] * b[244] + a[253] * b[264] + a[254] * b[284] + a[255] * b[304] + a[256] * b[324] + a[257] * b[344] + a[258] * b[364] + a[259] * b[384];
                    c[245] <= a[240] * b[5] + a[241] * b[25] + a[242] * b[45] + a[243] * b[65] + a[244] * b[85] + a[245] * b[105] + a[246] * b[125] + a[247] * b[145] + a[248] * b[165] + a[249] * b[185] + a[250] * b[205] + a[251] * b[225] + a[252] * b[245] + a[253] * b[265] + a[254] * b[285] + a[255] * b[305] + a[256] * b[325] + a[257] * b[345] + a[258] * b[365] + a[259] * b[385];
                    c[246] <= a[240] * b[6] + a[241] * b[26] + a[242] * b[46] + a[243] * b[66] + a[244] * b[86] + a[245] * b[106] + a[246] * b[126] + a[247] * b[146] + a[248] * b[166] + a[249] * b[186] + a[250] * b[206] + a[251] * b[226] + a[252] * b[246] + a[253] * b[266] + a[254] * b[286] + a[255] * b[306] + a[256] * b[326] + a[257] * b[346] + a[258] * b[366] + a[259] * b[386];
                    c[247] <= a[240] * b[7] + a[241] * b[27] + a[242] * b[47] + a[243] * b[67] + a[244] * b[87] + a[245] * b[107] + a[246] * b[127] + a[247] * b[147] + a[248] * b[167] + a[249] * b[187] + a[250] * b[207] + a[251] * b[227] + a[252] * b[247] + a[253] * b[267] + a[254] * b[287] + a[255] * b[307] + a[256] * b[327] + a[257] * b[347] + a[258] * b[367] + a[259] * b[387];
                    c[248] <= a[240] * b[8] + a[241] * b[28] + a[242] * b[48] + a[243] * b[68] + a[244] * b[88] + a[245] * b[108] + a[246] * b[128] + a[247] * b[148] + a[248] * b[168] + a[249] * b[188] + a[250] * b[208] + a[251] * b[228] + a[252] * b[248] + a[253] * b[268] + a[254] * b[288] + a[255] * b[308] + a[256] * b[328] + a[257] * b[348] + a[258] * b[368] + a[259] * b[388];
                    c[249] <= a[240] * b[9] + a[241] * b[29] + a[242] * b[49] + a[243] * b[69] + a[244] * b[89] + a[245] * b[109] + a[246] * b[129] + a[247] * b[149] + a[248] * b[169] + a[249] * b[189] + a[250] * b[209] + a[251] * b[229] + a[252] * b[249] + a[253] * b[269] + a[254] * b[289] + a[255] * b[309] + a[256] * b[329] + a[257] * b[349] + a[258] * b[369] + a[259] * b[389];
                    c[250] <= a[240] * b[10] + a[241] * b[30] + a[242] * b[50] + a[243] * b[70] + a[244] * b[90] + a[245] * b[110] + a[246] * b[130] + a[247] * b[150] + a[248] * b[170] + a[249] * b[190] + a[250] * b[210] + a[251] * b[230] + a[252] * b[250] + a[253] * b[270] + a[254] * b[290] + a[255] * b[310] + a[256] * b[330] + a[257] * b[350] + a[258] * b[370] + a[259] * b[390];
                    c[251] <= a[240] * b[11] + a[241] * b[31] + a[242] * b[51] + a[243] * b[71] + a[244] * b[91] + a[245] * b[111] + a[246] * b[131] + a[247] * b[151] + a[248] * b[171] + a[249] * b[191] + a[250] * b[211] + a[251] * b[231] + a[252] * b[251] + a[253] * b[271] + a[254] * b[291] + a[255] * b[311] + a[256] * b[331] + a[257] * b[351] + a[258] * b[371] + a[259] * b[391];
                    c[252] <= a[240] * b[12] + a[241] * b[32] + a[242] * b[52] + a[243] * b[72] + a[244] * b[92] + a[245] * b[112] + a[246] * b[132] + a[247] * b[152] + a[248] * b[172] + a[249] * b[192] + a[250] * b[212] + a[251] * b[232] + a[252] * b[252] + a[253] * b[272] + a[254] * b[292] + a[255] * b[312] + a[256] * b[332] + a[257] * b[352] + a[258] * b[372] + a[259] * b[392];
                    c[253] <= a[240] * b[13] + a[241] * b[33] + a[242] * b[53] + a[243] * b[73] + a[244] * b[93] + a[245] * b[113] + a[246] * b[133] + a[247] * b[153] + a[248] * b[173] + a[249] * b[193] + a[250] * b[213] + a[251] * b[233] + a[252] * b[253] + a[253] * b[273] + a[254] * b[293] + a[255] * b[313] + a[256] * b[333] + a[257] * b[353] + a[258] * b[373] + a[259] * b[393];
                    c[254] <= a[240] * b[14] + a[241] * b[34] + a[242] * b[54] + a[243] * b[74] + a[244] * b[94] + a[245] * b[114] + a[246] * b[134] + a[247] * b[154] + a[248] * b[174] + a[249] * b[194] + a[250] * b[214] + a[251] * b[234] + a[252] * b[254] + a[253] * b[274] + a[254] * b[294] + a[255] * b[314] + a[256] * b[334] + a[257] * b[354] + a[258] * b[374] + a[259] * b[394];
                    c[255] <= a[240] * b[15] + a[241] * b[35] + a[242] * b[55] + a[243] * b[75] + a[244] * b[95] + a[245] * b[115] + a[246] * b[135] + a[247] * b[155] + a[248] * b[175] + a[249] * b[195] + a[250] * b[215] + a[251] * b[235] + a[252] * b[255] + a[253] * b[275] + a[254] * b[295] + a[255] * b[315] + a[256] * b[335] + a[257] * b[355] + a[258] * b[375] + a[259] * b[395];
                    c[256] <= a[240] * b[16] + a[241] * b[36] + a[242] * b[56] + a[243] * b[76] + a[244] * b[96] + a[245] * b[116] + a[246] * b[136] + a[247] * b[156] + a[248] * b[176] + a[249] * b[196] + a[250] * b[216] + a[251] * b[236] + a[252] * b[256] + a[253] * b[276] + a[254] * b[296] + a[255] * b[316] + a[256] * b[336] + a[257] * b[356] + a[258] * b[376] + a[259] * b[396];
                    c[257] <= a[240] * b[17] + a[241] * b[37] + a[242] * b[57] + a[243] * b[77] + a[244] * b[97] + a[245] * b[117] + a[246] * b[137] + a[247] * b[157] + a[248] * b[177] + a[249] * b[197] + a[250] * b[217] + a[251] * b[237] + a[252] * b[257] + a[253] * b[277] + a[254] * b[297] + a[255] * b[317] + a[256] * b[337] + a[257] * b[357] + a[258] * b[377] + a[259] * b[397];
                    c[258] <= a[240] * b[18] + a[241] * b[38] + a[242] * b[58] + a[243] * b[78] + a[244] * b[98] + a[245] * b[118] + a[246] * b[138] + a[247] * b[158] + a[248] * b[178] + a[249] * b[198] + a[250] * b[218] + a[251] * b[238] + a[252] * b[258] + a[253] * b[278] + a[254] * b[298] + a[255] * b[318] + a[256] * b[338] + a[257] * b[358] + a[258] * b[378] + a[259] * b[398];
                    c[259] <= a[240] * b[19] + a[241] * b[39] + a[242] * b[59] + a[243] * b[79] + a[244] * b[99] + a[245] * b[119] + a[246] * b[139] + a[247] * b[159] + a[248] * b[179] + a[249] * b[199] + a[250] * b[219] + a[251] * b[239] + a[252] * b[259] + a[253] * b[279] + a[254] * b[299] + a[255] * b[319] + a[256] * b[339] + a[257] * b[359] + a[258] * b[379] + a[259] * b[399];
                    c[260] <= a[260] * b[0] + a[261] * b[20] + a[262] * b[40] + a[263] * b[60] + a[264] * b[80] + a[265] * b[100] + a[266] * b[120] + a[267] * b[140] + a[268] * b[160] + a[269] * b[180] + a[270] * b[200] + a[271] * b[220] + a[272] * b[240] + a[273] * b[260] + a[274] * b[280] + a[275] * b[300] + a[276] * b[320] + a[277] * b[340] + a[278] * b[360] + a[279] * b[380];
                    c[261] <= a[260] * b[1] + a[261] * b[21] + a[262] * b[41] + a[263] * b[61] + a[264] * b[81] + a[265] * b[101] + a[266] * b[121] + a[267] * b[141] + a[268] * b[161] + a[269] * b[181] + a[270] * b[201] + a[271] * b[221] + a[272] * b[241] + a[273] * b[261] + a[274] * b[281] + a[275] * b[301] + a[276] * b[321] + a[277] * b[341] + a[278] * b[361] + a[279] * b[381];
                    c[262] <= a[260] * b[2] + a[261] * b[22] + a[262] * b[42] + a[263] * b[62] + a[264] * b[82] + a[265] * b[102] + a[266] * b[122] + a[267] * b[142] + a[268] * b[162] + a[269] * b[182] + a[270] * b[202] + a[271] * b[222] + a[272] * b[242] + a[273] * b[262] + a[274] * b[282] + a[275] * b[302] + a[276] * b[322] + a[277] * b[342] + a[278] * b[362] + a[279] * b[382];
                    c[263] <= a[260] * b[3] + a[261] * b[23] + a[262] * b[43] + a[263] * b[63] + a[264] * b[83] + a[265] * b[103] + a[266] * b[123] + a[267] * b[143] + a[268] * b[163] + a[269] * b[183] + a[270] * b[203] + a[271] * b[223] + a[272] * b[243] + a[273] * b[263] + a[274] * b[283] + a[275] * b[303] + a[276] * b[323] + a[277] * b[343] + a[278] * b[363] + a[279] * b[383];
                    c[264] <= a[260] * b[4] + a[261] * b[24] + a[262] * b[44] + a[263] * b[64] + a[264] * b[84] + a[265] * b[104] + a[266] * b[124] + a[267] * b[144] + a[268] * b[164] + a[269] * b[184] + a[270] * b[204] + a[271] * b[224] + a[272] * b[244] + a[273] * b[264] + a[274] * b[284] + a[275] * b[304] + a[276] * b[324] + a[277] * b[344] + a[278] * b[364] + a[279] * b[384];
                    c[265] <= a[260] * b[5] + a[261] * b[25] + a[262] * b[45] + a[263] * b[65] + a[264] * b[85] + a[265] * b[105] + a[266] * b[125] + a[267] * b[145] + a[268] * b[165] + a[269] * b[185] + a[270] * b[205] + a[271] * b[225] + a[272] * b[245] + a[273] * b[265] + a[274] * b[285] + a[275] * b[305] + a[276] * b[325] + a[277] * b[345] + a[278] * b[365] + a[279] * b[385];
                    c[266] <= a[260] * b[6] + a[261] * b[26] + a[262] * b[46] + a[263] * b[66] + a[264] * b[86] + a[265] * b[106] + a[266] * b[126] + a[267] * b[146] + a[268] * b[166] + a[269] * b[186] + a[270] * b[206] + a[271] * b[226] + a[272] * b[246] + a[273] * b[266] + a[274] * b[286] + a[275] * b[306] + a[276] * b[326] + a[277] * b[346] + a[278] * b[366] + a[279] * b[386];
                    c[267] <= a[260] * b[7] + a[261] * b[27] + a[262] * b[47] + a[263] * b[67] + a[264] * b[87] + a[265] * b[107] + a[266] * b[127] + a[267] * b[147] + a[268] * b[167] + a[269] * b[187] + a[270] * b[207] + a[271] * b[227] + a[272] * b[247] + a[273] * b[267] + a[274] * b[287] + a[275] * b[307] + a[276] * b[327] + a[277] * b[347] + a[278] * b[367] + a[279] * b[387];
                    c[268] <= a[260] * b[8] + a[261] * b[28] + a[262] * b[48] + a[263] * b[68] + a[264] * b[88] + a[265] * b[108] + a[266] * b[128] + a[267] * b[148] + a[268] * b[168] + a[269] * b[188] + a[270] * b[208] + a[271] * b[228] + a[272] * b[248] + a[273] * b[268] + a[274] * b[288] + a[275] * b[308] + a[276] * b[328] + a[277] * b[348] + a[278] * b[368] + a[279] * b[388];
                    c[269] <= a[260] * b[9] + a[261] * b[29] + a[262] * b[49] + a[263] * b[69] + a[264] * b[89] + a[265] * b[109] + a[266] * b[129] + a[267] * b[149] + a[268] * b[169] + a[269] * b[189] + a[270] * b[209] + a[271] * b[229] + a[272] * b[249] + a[273] * b[269] + a[274] * b[289] + a[275] * b[309] + a[276] * b[329] + a[277] * b[349] + a[278] * b[369] + a[279] * b[389];
                    c[270] <= a[260] * b[10] + a[261] * b[30] + a[262] * b[50] + a[263] * b[70] + a[264] * b[90] + a[265] * b[110] + a[266] * b[130] + a[267] * b[150] + a[268] * b[170] + a[269] * b[190] + a[270] * b[210] + a[271] * b[230] + a[272] * b[250] + a[273] * b[270] + a[274] * b[290] + a[275] * b[310] + a[276] * b[330] + a[277] * b[350] + a[278] * b[370] + a[279] * b[390];
                    c[271] <= a[260] * b[11] + a[261] * b[31] + a[262] * b[51] + a[263] * b[71] + a[264] * b[91] + a[265] * b[111] + a[266] * b[131] + a[267] * b[151] + a[268] * b[171] + a[269] * b[191] + a[270] * b[211] + a[271] * b[231] + a[272] * b[251] + a[273] * b[271] + a[274] * b[291] + a[275] * b[311] + a[276] * b[331] + a[277] * b[351] + a[278] * b[371] + a[279] * b[391];
                    c[272] <= a[260] * b[12] + a[261] * b[32] + a[262] * b[52] + a[263] * b[72] + a[264] * b[92] + a[265] * b[112] + a[266] * b[132] + a[267] * b[152] + a[268] * b[172] + a[269] * b[192] + a[270] * b[212] + a[271] * b[232] + a[272] * b[252] + a[273] * b[272] + a[274] * b[292] + a[275] * b[312] + a[276] * b[332] + a[277] * b[352] + a[278] * b[372] + a[279] * b[392];
                    c[273] <= a[260] * b[13] + a[261] * b[33] + a[262] * b[53] + a[263] * b[73] + a[264] * b[93] + a[265] * b[113] + a[266] * b[133] + a[267] * b[153] + a[268] * b[173] + a[269] * b[193] + a[270] * b[213] + a[271] * b[233] + a[272] * b[253] + a[273] * b[273] + a[274] * b[293] + a[275] * b[313] + a[276] * b[333] + a[277] * b[353] + a[278] * b[373] + a[279] * b[393];
                    c[274] <= a[260] * b[14] + a[261] * b[34] + a[262] * b[54] + a[263] * b[74] + a[264] * b[94] + a[265] * b[114] + a[266] * b[134] + a[267] * b[154] + a[268] * b[174] + a[269] * b[194] + a[270] * b[214] + a[271] * b[234] + a[272] * b[254] + a[273] * b[274] + a[274] * b[294] + a[275] * b[314] + a[276] * b[334] + a[277] * b[354] + a[278] * b[374] + a[279] * b[394];
                    c[275] <= a[260] * b[15] + a[261] * b[35] + a[262] * b[55] + a[263] * b[75] + a[264] * b[95] + a[265] * b[115] + a[266] * b[135] + a[267] * b[155] + a[268] * b[175] + a[269] * b[195] + a[270] * b[215] + a[271] * b[235] + a[272] * b[255] + a[273] * b[275] + a[274] * b[295] + a[275] * b[315] + a[276] * b[335] + a[277] * b[355] + a[278] * b[375] + a[279] * b[395];
                    c[276] <= a[260] * b[16] + a[261] * b[36] + a[262] * b[56] + a[263] * b[76] + a[264] * b[96] + a[265] * b[116] + a[266] * b[136] + a[267] * b[156] + a[268] * b[176] + a[269] * b[196] + a[270] * b[216] + a[271] * b[236] + a[272] * b[256] + a[273] * b[276] + a[274] * b[296] + a[275] * b[316] + a[276] * b[336] + a[277] * b[356] + a[278] * b[376] + a[279] * b[396];
                    c[277] <= a[260] * b[17] + a[261] * b[37] + a[262] * b[57] + a[263] * b[77] + a[264] * b[97] + a[265] * b[117] + a[266] * b[137] + a[267] * b[157] + a[268] * b[177] + a[269] * b[197] + a[270] * b[217] + a[271] * b[237] + a[272] * b[257] + a[273] * b[277] + a[274] * b[297] + a[275] * b[317] + a[276] * b[337] + a[277] * b[357] + a[278] * b[377] + a[279] * b[397];
                    c[278] <= a[260] * b[18] + a[261] * b[38] + a[262] * b[58] + a[263] * b[78] + a[264] * b[98] + a[265] * b[118] + a[266] * b[138] + a[267] * b[158] + a[268] * b[178] + a[269] * b[198] + a[270] * b[218] + a[271] * b[238] + a[272] * b[258] + a[273] * b[278] + a[274] * b[298] + a[275] * b[318] + a[276] * b[338] + a[277] * b[358] + a[278] * b[378] + a[279] * b[398];
                    c[279] <= a[260] * b[19] + a[261] * b[39] + a[262] * b[59] + a[263] * b[79] + a[264] * b[99] + a[265] * b[119] + a[266] * b[139] + a[267] * b[159] + a[268] * b[179] + a[269] * b[199] + a[270] * b[219] + a[271] * b[239] + a[272] * b[259] + a[273] * b[279] + a[274] * b[299] + a[275] * b[319] + a[276] * b[339] + a[277] * b[359] + a[278] * b[379] + a[279] * b[399];
                end
            endcase
        end
    end

    always @(posedge clk) begin
        if (rst) begin
            state <= 0;
        end else begin
            case (state)
                fin: begin
                    if (matmult_accept) begin
                        state <= idle;
                    end
                end
                idle: begin
                    if (matmult_ready) begin
                        state <= calc;
                    end
                end
                calc: begin
                    state <= fin;
                end
            endcase
        end
    end

endmodule
